module __sha256__main(
  input wire [511:0] message,
  output wire [255:0] out
);
  wire [28:0] add_56574;
  wire [30:0] add_56578;
  wire [31:0] e__66;
  wire [31:0] f__1;
  wire [5:0] S1__67;
  wire [4:0] S1__66;
  wire [13:0] S1__65;
  wire [6:0] S1__64;
  wire [31:0] S1__1;
  wire [31:0] ch__1;
  wire [29:0] add_56608;
  wire [31:0] temp1__336;
  wire [31:0] temp1__337;
  wire [31:0] temp1__338;
  wire [30:0] add_56615;
  wire [31:0] e__67;
  wire [5:0] S1__71;
  wire [4:0] S1__70;
  wire [13:0] S1__69;
  wire [6:0] S1__68;
  wire [31:0] S1__2;
  wire [31:0] ch__2;
  wire [31:0] w_im15__1;
  wire [31:0] temp1__331;
  wire [31:0] temp1__332;
  wire [31:0] temp1__333;
  wire [31:0] temp1__334;
  wire [31:0] c__67;
  wire [31:0] e__68;
  wire [5:0] S1__75;
  wire [4:0] S1__74;
  wire [13:0] S1__73;
  wire [6:0] S1__72;
  wire [31:0] S1__3;
  wire [31:0] ch__3;
  wire [29:0] add_56676;
  wire [31:0] temp1__328;
  wire [31:0] temp1__329;
  wire [31:0] temp1__330;
  wire [31:0] b__67;
  wire [31:0] e__69;
  wire [5:0] S1__79;
  wire [4:0] S1__78;
  wire [13:0] S1__77;
  wire [6:0] S1__76;
  wire [31:0] S1__4;
  wire [31:0] temp1__17;
  wire [31:0] ch__4;
  wire [31:0] w_im15__3;
  wire [31:0] temp1__323;
  wire [31:0] temp2;
  wire [31:0] temp1__18;
  wire [31:0] temp1__262;
  wire [31:0] a__1;
  wire [31:0] temp1__20;
  wire [31:0] e__5;
  wire [31:0] b__1;
  wire [31:0] c__1;
  wire [5:0] S1__83;
  wire [4:0] S1__82;
  wire [13:0] S1__81;
  wire [6:0] S1__80;
  wire [1:0] S0__67;
  wire [10:0] S0__66;
  wire [8:0] S0__65;
  wire [9:0] S0__64;
  wire [31:0] and_56752;
  wire [31:0] S1__5;
  wire [31:0] S0__1;
  wire [31:0] maj__1;
  wire [31:0] temp1__21;
  wire [31:0] ch__5;
  wire [31:0] w_im15__4;
  wire [31:0] temp2__1;
  wire [31:0] temp1__22;
  wire [31:0] temp1__263;
  wire [31:0] a__2;
  wire [31:0] temp1__24;
  wire [31:0] e__6;
  wire [31:0] b__66;
  wire [1:0] S0__71;
  wire [10:0] S0__70;
  wire [8:0] S0__69;
  wire [9:0] S0__68;
  wire [31:0] and_56802;
  wire [5:0] S1__87;
  wire [4:0] S1__86;
  wire [13:0] S1__85;
  wire [6:0] S1__84;
  wire [29:0] add_56810;
  wire [31:0] S0__2;
  wire [31:0] maj__2;
  wire [31:0] S1__6;
  wire [31:0] ch__6;
  wire [31:0] temp1__264;
  wire [31:0] temp2__2;
  wire [31:0] temp1__437;
  wire [31:0] temp1__438;
  wire [31:0] a__3;
  wire [31:0] temp1__439;
  wire [31:0] e__7;
  wire [5:0] S1__91;
  wire [4:0] S1__90;
  wire [13:0] S1__89;
  wire [6:0] S1__88;
  wire [1:0] S0__75;
  wire [10:0] S0__74;
  wire [8:0] S0__73;
  wire [9:0] S0__72;
  wire [31:0] and_56856;
  wire [31:0] S1__7;
  wire [31:0] S0__3;
  wire [31:0] maj__3;
  wire [31:0] temp1__29;
  wire [31:0] ch__7;
  wire [31:0] w_im15__6;
  wire [31:0] temp2__3;
  wire [31:0] temp1__30;
  wire [31:0] temp1__265;
  wire [31:0] a__4;
  wire [31:0] temp1__32;
  wire [31:0] e__8;
  wire [1:0] S0__79;
  wire [10:0] S0__78;
  wire [8:0] S0__77;
  wire [9:0] S0__76;
  wire [31:0] and_56904;
  wire [5:0] S1__95;
  wire [4:0] S1__94;
  wire [13:0] S1__93;
  wire [6:0] S1__92;
  wire [28:0] add_56912;
  wire [31:0] S0__4;
  wire [31:0] maj__4;
  wire [31:0] S1__8;
  wire [31:0] ch__8;
  wire [31:0] temp1__266;
  wire [31:0] temp2__4;
  wire [31:0] temp1__434;
  wire [31:0] temp1__435;
  wire [31:0] a__5;
  wire [31:0] temp1__436;
  wire [31:0] e__9;
  wire [5:0] S1__99;
  wire [4:0] S1__98;
  wire [13:0] S1__97;
  wire [6:0] S1__96;
  wire [1:0] S0__83;
  wire [10:0] S0__82;
  wire [8:0] S0__81;
  wire [9:0] S0__80;
  wire [31:0] and_56958;
  wire [31:0] S1__9;
  wire [31:0] S0__5;
  wire [31:0] maj__5;
  wire [31:0] temp1__37;
  wire [31:0] ch__9;
  wire [31:0] w_im15__8;
  wire [31:0] temp2__5;
  wire [31:0] temp1__38;
  wire [31:0] temp1__267;
  wire [31:0] a__6;
  wire [31:0] temp1__40;
  wire [31:0] e__10;
  wire [1:0] S0__87;
  wire [10:0] S0__86;
  wire [8:0] S0__85;
  wire [9:0] S0__84;
  wire [31:0] and_57006;
  wire [5:0] S1__103;
  wire [4:0] S1__102;
  wire [13:0] S1__101;
  wire [6:0] S1__100;
  wire [30:0] add_57014;
  wire [31:0] S0__6;
  wire [31:0] maj__6;
  wire [31:0] S1__10;
  wire [31:0] ch__10;
  wire [31:0] temp1__268;
  wire [31:0] temp2__6;
  wire [31:0] temp1__431;
  wire [31:0] temp1__432;
  wire [31:0] a__7;
  wire [31:0] temp1__433;
  wire [31:0] e__11;
  wire [5:0] S1__107;
  wire [4:0] S1__106;
  wire [13:0] S1__105;
  wire [6:0] S1__104;
  wire [1:0] S0__91;
  wire [10:0] S0__90;
  wire [8:0] S0__89;
  wire [9:0] S0__88;
  wire [31:0] and_57060;
  wire [31:0] S1__11;
  wire [31:0] S0__7;
  wire [31:0] maj__7;
  wire [31:0] temp1__45;
  wire [31:0] ch__11;
  wire [31:0] w_im15__10;
  wire [31:0] temp2__7;
  wire [31:0] temp1__46;
  wire [31:0] temp1__269;
  wire [31:0] a__8;
  wire [31:0] temp1__48;
  wire [31:0] e__12;
  wire [1:0] S0__95;
  wire [10:0] S0__94;
  wire [8:0] S0__93;
  wire [9:0] S0__92;
  wire [31:0] and_57108;
  wire [5:0] S1__111;
  wire [4:0] S1__110;
  wire [13:0] S1__109;
  wire [6:0] S1__108;
  wire [29:0] add_57116;
  wire [31:0] S0__8;
  wire [31:0] maj__8;
  wire [31:0] S1__12;
  wire [31:0] ch__12;
  wire [31:0] temp1__270;
  wire [31:0] temp2__8;
  wire [31:0] temp1__428;
  wire [31:0] temp1__429;
  wire [31:0] a__9;
  wire [31:0] temp1__430;
  wire [31:0] e__13;
  wire [1:0] S0__99;
  wire [10:0] S0__98;
  wire [8:0] S0__97;
  wire [9:0] S0__96;
  wire [31:0] and_57160;
  wire [5:0] S1__115;
  wire [4:0] S1__114;
  wire [13:0] S1__113;
  wire [6:0] S1__112;
  wire [30:0] add_57168;
  wire [31:0] S0__9;
  wire [31:0] maj__9;
  wire [31:0] S1__13;
  wire [31:0] ch__13;
  wire [31:0] temp1__271;
  wire [31:0] temp2__9;
  wire [31:0] temp1__425;
  wire [31:0] temp1__426;
  wire [31:0] a__10;
  wire [31:0] temp1__427;
  wire [31:0] e__14;
  wire [5:0] S1__119;
  wire [4:0] S1__118;
  wire [13:0] S1__117;
  wire [6:0] S1__116;
  wire [1:0] S0__103;
  wire [10:0] S0__102;
  wire [8:0] S0__101;
  wire [9:0] S0__100;
  wire [31:0] and_57214;
  wire [31:0] S1__14;
  wire [31:0] S0__10;
  wire [31:0] maj__10;
  wire [31:0] temp1__57;
  wire [31:0] ch__14;
  wire [31:0] w_init_im2;
  wire [31:0] temp2__10;
  wire [31:0] temp1__58;
  wire [31:0] temp1__272;
  wire [31:0] a__11;
  wire [31:0] temp1__60;
  wire [31:0] e__15;
  wire [1:0] S0__107;
  wire [10:0] S0__106;
  wire [8:0] S0__105;
  wire [9:0] S0__104;
  wire [31:0] and_57262;
  wire [5:0] S1__123;
  wire [4:0] S1__122;
  wire [13:0] S1__121;
  wire [6:0] S1__120;
  wire [29:0] add_57270;
  wire [31:0] S0__11;
  wire [31:0] maj__11;
  wire [31:0] S1__15;
  wire [31:0] ch__15;
  wire [31:0] temp1__273;
  wire [31:0] temp2__11;
  wire [31:0] temp1__422;
  wire [31:0] temp1__423;
  wire [31:0] a__12;
  wire [31:0] temp1__424;
  wire [31:0] e__16;
  wire [2:0] s_0__51;
  wire [3:0] s_0__50;
  wire [10:0] s_0__49;
  wire [13:0] s_0__48;
  wire [9:0] s_1__51;
  wire [6:0] s_1__50;
  wire [1:0] s_1__49;
  wire [12:0] s_1__48;
  wire [5:0] S1__127;
  wire [4:0] S1__126;
  wire [13:0] S1__125;
  wire [6:0] S1__124;
  wire [31:0] s_0__1;
  wire [31:0] s_1__1;
  wire [1:0] S0__111;
  wire [10:0] S0__110;
  wire [8:0] S0__109;
  wire [9:0] S0__108;
  wire [31:0] and_57349;
  wire [31:0] S1__16;
  wire [31:0] value__1;
  wire [31:0] value__2;
  wire [31:0] S0__12;
  wire [31:0] maj__12;
  wire [31:0] temp1__65;
  wire [31:0] ch__16;
  wire [31:0] value__3;
  wire [2:0] s_0__55;
  wire [3:0] s_0__54;
  wire [10:0] s_0__53;
  wire [13:0] s_0__52;
  wire [9:0] s_1__55;
  wire [6:0] s_1__54;
  wire [1:0] s_1__53;
  wire [12:0] s_1__52;
  wire [31:0] temp2__12;
  wire [31:0] temp1__66;
  wire [31:0] temp1__274;
  wire [31:0] w_init_im15;
  wire [31:0] s_0__2;
  wire [31:0] w_im15__9;
  wire [31:0] s_1__2;
  wire [31:0] a__13;
  wire [31:0] temp1__68;
  wire [31:0] value__4;
  wire [31:0] value__5;
  wire [31:0] e__17;
  wire [31:0] value__6;
  wire [1:0] S0__115;
  wire [10:0] S0__114;
  wire [8:0] S0__113;
  wire [9:0] S0__112;
  wire [31:0] and_57435;
  wire [5:0] S1__131;
  wire [4:0] S1__130;
  wire [13:0] S1__129;
  wire [6:0] S1__128;
  wire [30:0] add_57443;
  wire [31:0] S0__13;
  wire [31:0] maj__13;
  wire [31:0] S1__17;
  wire [31:0] ch__17;
  wire [31:0] temp1__275;
  wire [2:0] s_0__59;
  wire [3:0] s_0__58;
  wire [10:0] s_0__57;
  wire [13:0] s_0__56;
  wire [9:0] s_1__59;
  wire [6:0] s_1__58;
  wire [1:0] s_1__57;
  wire [12:0] s_1__56;
  wire [31:0] temp2__13;
  wire [31:0] temp1__419;
  wire [31:0] temp1__420;
  wire [31:0] s_0__3;
  wire [31:0] s_1__3;
  wire [31:0] a__14;
  wire [31:0] temp1__421;
  wire [31:0] value__7;
  wire [31:0] value__8;
  wire [31:0] e__18;
  wire [31:0] value__9;
  wire [1:0] S0__119;
  wire [10:0] S0__118;
  wire [8:0] S0__117;
  wire [9:0] S0__116;
  wire [31:0] and_57522;
  wire [5:0] S1__135;
  wire [4:0] S1__134;
  wire [13:0] S1__133;
  wire [6:0] S1__132;
  wire [30:0] add_57530;
  wire [31:0] S0__14;
  wire [31:0] maj__14;
  wire [31:0] S1__18;
  wire [31:0] ch__18;
  wire [31:0] temp1__276;
  wire [2:0] s_0__63;
  wire [3:0] s_0__62;
  wire [10:0] s_0__61;
  wire [13:0] s_0__60;
  wire [9:0] s_1__63;
  wire [6:0] s_1__62;
  wire [1:0] s_1__61;
  wire [12:0] s_1__60;
  wire [31:0] temp2__14;
  wire [31:0] temp1__416;
  wire [31:0] temp1__417;
  wire [31:0] w_im15__2;
  wire [31:0] s_0__4;
  wire [31:0] w_im15__11;
  wire [31:0] s_1__4;
  wire [31:0] a__15;
  wire [31:0] temp1__418;
  wire [31:0] value__10;
  wire [31:0] value__11;
  wire [31:0] e__19;
  wire [31:0] value__12;
  wire [1:0] S0__123;
  wire [10:0] S0__122;
  wire [8:0] S0__121;
  wire [9:0] S0__120;
  wire [31:0] and_57611;
  wire [5:0] S1__139;
  wire [4:0] S1__138;
  wire [13:0] S1__137;
  wire [6:0] S1__136;
  wire [29:0] add_57619;
  wire [31:0] S0__15;
  wire [31:0] maj__15;
  wire [31:0] S1__19;
  wire [31:0] ch__19;
  wire [31:0] temp1__277;
  wire [31:0] temp2__15;
  wire [31:0] temp1__413;
  wire [31:0] temp1__414;
  wire [31:0] a__16;
  wire [31:0] temp1__415;
  wire [31:0] e__20;
  wire [2:0] s_0__67;
  wire [3:0] s_0__66;
  wire [10:0] s_0__65;
  wire [13:0] s_0__64;
  wire [9:0] s_1__67;
  wire [6:0] s_1__66;
  wire [1:0] s_1__65;
  wire [12:0] s_1__64;
  wire [5:0] S1__143;
  wire [4:0] S1__142;
  wire [13:0] S1__141;
  wire [6:0] S1__140;
  wire [31:0] s_0__5;
  wire [31:0] w_im15__12;
  wire [31:0] s_1__5;
  wire [1:0] S0__127;
  wire [10:0] S0__126;
  wire [8:0] S0__125;
  wire [9:0] S0__124;
  wire [31:0] and_57698;
  wire [31:0] S1__20;
  wire [31:0] value__13;
  wire [31:0] value__14;
  wire [31:0] S0__16;
  wire [31:0] maj__16;
  wire [31:0] temp1__81;
  wire [31:0] ch__20;
  wire [31:0] value__15;
  wire [2:0] s_0__71;
  wire [3:0] s_0__70;
  wire [10:0] s_0__69;
  wire [13:0] s_0__68;
  wire [9:0] s_1__71;
  wire [6:0] s_1__70;
  wire [1:0] s_1__69;
  wire [12:0] s_1__68;
  wire [31:0] temp2__16;
  wire [31:0] temp1__82;
  wire [31:0] temp1__278;
  wire [31:0] s_0__6;
  wire [31:0] s_1__6;
  wire [31:0] a__17;
  wire [31:0] temp1__84;
  wire [31:0] value__16;
  wire [31:0] value__17;
  wire [31:0] e__21;
  wire [31:0] value__18;
  wire [1:0] S0__131;
  wire [10:0] S0__130;
  wire [8:0] S0__129;
  wire [9:0] S0__128;
  wire [31:0] and_57782;
  wire [5:0] S1__147;
  wire [4:0] S1__146;
  wire [13:0] S1__145;
  wire [6:0] S1__144;
  wire [30:0] add_57790;
  wire [31:0] S0__17;
  wire [31:0] maj__17;
  wire [31:0] S1__21;
  wire [31:0] ch__21;
  wire [31:0] temp1__279;
  wire [2:0] s_0__75;
  wire [3:0] s_0__74;
  wire [10:0] s_0__73;
  wire [13:0] s_0__72;
  wire [9:0] s_1__75;
  wire [6:0] s_1__74;
  wire [1:0] s_1__73;
  wire [12:0] s_1__72;
  wire [31:0] temp2__17;
  wire [31:0] temp1__410;
  wire [31:0] temp1__411;
  wire [31:0] w_im15__5;
  wire [31:0] s_0__7;
  wire [31:0] w_im2__1;
  wire [31:0] s_1__7;
  wire [31:0] a__18;
  wire [31:0] temp1__412;
  wire [31:0] value__19;
  wire [31:0] value__20;
  wire [31:0] e__22;
  wire [31:0] value__21;
  wire [1:0] S0__135;
  wire [10:0] S0__134;
  wire [8:0] S0__133;
  wire [9:0] S0__132;
  wire [31:0] and_57871;
  wire [5:0] S1__151;
  wire [4:0] S1__150;
  wire [13:0] S1__149;
  wire [6:0] S1__148;
  wire [29:0] add_57879;
  wire [31:0] S0__18;
  wire [31:0] maj__18;
  wire [31:0] S1__22;
  wire [31:0] ch__22;
  wire [31:0] temp1__280;
  wire [2:0] s_0__79;
  wire [3:0] s_0__78;
  wire [10:0] s_0__77;
  wire [13:0] s_0__76;
  wire [9:0] s_1__79;
  wire [6:0] s_1__78;
  wire [1:0] s_1__77;
  wire [12:0] s_1__76;
  wire [31:0] temp2__18;
  wire [31:0] temp1__407;
  wire [31:0] temp1__408;
  wire [31:0] s_0__8;
  wire [31:0] s_1__8;
  wire [31:0] a__19;
  wire [31:0] temp1__409;
  wire [31:0] value__22;
  wire [31:0] value__23;
  wire [31:0] e__23;
  wire [31:0] value__24;
  wire [1:0] S0__139;
  wire [10:0] S0__138;
  wire [8:0] S0__137;
  wire [9:0] S0__136;
  wire [31:0] and_57958;
  wire [5:0] S1__155;
  wire [4:0] S1__154;
  wire [13:0] S1__153;
  wire [6:0] S1__152;
  wire [30:0] add_57966;
  wire [31:0] S0__19;
  wire [31:0] maj__19;
  wire [31:0] S1__23;
  wire [31:0] ch__23;
  wire [31:0] temp1__281;
  wire [2:0] s_0__83;
  wire [3:0] s_0__82;
  wire [10:0] s_0__81;
  wire [13:0] s_0__80;
  wire [9:0] s_1__83;
  wire [6:0] s_1__82;
  wire [1:0] s_1__81;
  wire [12:0] s_1__80;
  wire [31:0] temp2__19;
  wire [31:0] temp1__404;
  wire [31:0] temp1__405;
  wire [31:0] w_im15__7;
  wire [31:0] s_0__9;
  wire [31:0] s_1__9;
  wire [31:0] a__20;
  wire [31:0] temp1__406;
  wire [31:0] value__25;
  wire [31:0] value__26;
  wire [31:0] e__24;
  wire [31:0] value__27;
  wire [1:0] S0__143;
  wire [10:0] S0__142;
  wire [8:0] S0__141;
  wire [9:0] S0__140;
  wire [31:0] and_58045;
  wire [5:0] S1__159;
  wire [4:0] S1__158;
  wire [13:0] S1__157;
  wire [6:0] S1__156;
  wire [30:0] add_58053;
  wire [31:0] S0__20;
  wire [31:0] maj__20;
  wire [31:0] S1__24;
  wire [31:0] ch__24;
  wire [31:0] temp1__282;
  wire [31:0] temp2__20;
  wire [31:0] temp1__401;
  wire [31:0] temp1__402;
  wire [31:0] a__21;
  wire [31:0] temp1__403;
  wire [31:0] e__25;
  wire [2:0] s_0__87;
  wire [3:0] s_0__86;
  wire [10:0] s_0__85;
  wire [13:0] s_0__84;
  wire [9:0] s_1__87;
  wire [6:0] s_1__86;
  wire [1:0] s_1__85;
  wire [12:0] s_1__84;
  wire [5:0] S1__163;
  wire [4:0] S1__162;
  wire [13:0] S1__161;
  wire [6:0] S1__160;
  wire [31:0] s_0__10;
  wire [31:0] s_1__10;
  wire [1:0] S0__147;
  wire [10:0] S0__146;
  wire [8:0] S0__145;
  wire [9:0] S0__144;
  wire [31:0] and_58131;
  wire [31:0] S1__25;
  wire [31:0] value__28;
  wire [31:0] value__29;
  wire [31:0] S0__21;
  wire [31:0] maj__21;
  wire [31:0] temp1__101;
  wire [31:0] ch__25;
  wire [31:0] value__30;
  wire [2:0] s_0__91;
  wire [3:0] s_0__90;
  wire [10:0] s_0__89;
  wire [13:0] s_0__88;
  wire [9:0] s_1__91;
  wire [6:0] s_1__90;
  wire [1:0] s_1__89;
  wire [12:0] s_1__88;
  wire [31:0] temp2__21;
  wire [31:0] temp1__102;
  wire [31:0] temp1__283;
  wire [31:0] s_0__11;
  wire [31:0] s_1__11;
  wire [31:0] a__22;
  wire [31:0] temp1__104;
  wire [31:0] value__31;
  wire [31:0] value__32;
  wire [31:0] e__26;
  wire [31:0] value__33;
  wire [1:0] S0__151;
  wire [10:0] S0__150;
  wire [8:0] S0__149;
  wire [9:0] S0__148;
  wire [31:0] and_58216;
  wire [5:0] S1__167;
  wire [4:0] S1__166;
  wire [13:0] S1__165;
  wire [6:0] S1__164;
  wire [28:0] add_58224;
  wire [31:0] S0__22;
  wire [31:0] maj__22;
  wire [31:0] S1__26;
  wire [31:0] ch__26;
  wire [31:0] temp1__284;
  wire [31:0] temp2__22;
  wire [31:0] temp1__398;
  wire [31:0] temp1__399;
  wire [31:0] a__23;
  wire [31:0] temp1__400;
  wire [31:0] e__27;
  wire [2:0] s_0__95;
  wire [3:0] s_0__94;
  wire [10:0] s_0__93;
  wire [13:0] s_0__92;
  wire [9:0] s_1__95;
  wire [6:0] s_1__94;
  wire [1:0] s_1__93;
  wire [12:0] s_1__92;
  wire [5:0] S1__171;
  wire [4:0] S1__170;
  wire [13:0] S1__169;
  wire [6:0] S1__168;
  wire [31:0] s_0__12;
  wire [31:0] s_1__12;
  wire [1:0] S0__155;
  wire [10:0] S0__154;
  wire [8:0] S0__153;
  wire [9:0] S0__152;
  wire [31:0] and_58302;
  wire [31:0] S1__27;
  wire [31:0] value__34;
  wire [31:0] value__35;
  wire [31:0] S0__23;
  wire [31:0] maj__23;
  wire [31:0] temp1__109;
  wire [31:0] ch__27;
  wire [31:0] value__36;
  wire [31:0] temp2__23;
  wire [31:0] temp1__110;
  wire [31:0] temp1__285;
  wire [31:0] a__24;
  wire [31:0] temp1__112;
  wire [31:0] e__28;
  wire [2:0] s_0__99;
  wire [3:0] s_0__98;
  wire [10:0] s_0__97;
  wire [13:0] s_0__96;
  wire [9:0] s_1__99;
  wire [6:0] s_1__98;
  wire [1:0] s_1__97;
  wire [12:0] s_1__96;
  wire [5:0] S1__175;
  wire [4:0] S1__174;
  wire [13:0] S1__173;
  wire [6:0] S1__172;
  wire [31:0] s_0__13;
  wire [31:0] s_1__13;
  wire [1:0] S0__159;
  wire [10:0] S0__158;
  wire [8:0] S0__157;
  wire [9:0] S0__156;
  wire [31:0] and_58386;
  wire [31:0] S1__28;
  wire [31:0] value__37;
  wire [31:0] value__38;
  wire [31:0] S0__24;
  wire [31:0] maj__24;
  wire [31:0] temp1__113;
  wire [31:0] ch__28;
  wire [31:0] value__39;
  wire [31:0] temp2__24;
  wire [31:0] temp1__114;
  wire [31:0] temp1__286;
  wire [31:0] a__25;
  wire [31:0] temp1__116;
  wire [31:0] e__29;
  wire [2:0] s_0__103;
  wire [3:0] s_0__102;
  wire [10:0] s_0__101;
  wire [13:0] s_0__100;
  wire [9:0] s_1__103;
  wire [6:0] s_1__102;
  wire [1:0] s_1__101;
  wire [12:0] s_1__100;
  wire [5:0] S1__179;
  wire [4:0] S1__178;
  wire [13:0] S1__177;
  wire [6:0] S1__176;
  wire [31:0] s_0__14;
  wire [31:0] s_1__14;
  wire [1:0] S0__163;
  wire [10:0] S0__162;
  wire [8:0] S0__161;
  wire [9:0] S0__160;
  wire [31:0] and_58470;
  wire [31:0] S1__29;
  wire [31:0] value__40;
  wire [31:0] value__41;
  wire [31:0] S0__25;
  wire [31:0] maj__25;
  wire [31:0] temp1__117;
  wire [31:0] ch__29;
  wire [31:0] value__42;
  wire [31:0] temp2__25;
  wire [31:0] temp1__118;
  wire [31:0] temp1__287;
  wire [31:0] a__26;
  wire [31:0] temp1__120;
  wire [31:0] e__30;
  wire [2:0] s_0__107;
  wire [3:0] s_0__106;
  wire [10:0] s_0__105;
  wire [13:0] s_0__104;
  wire [9:0] s_1__107;
  wire [6:0] s_1__106;
  wire [1:0] s_1__105;
  wire [12:0] s_1__104;
  wire [5:0] S1__183;
  wire [4:0] S1__182;
  wire [13:0] S1__181;
  wire [6:0] S1__180;
  wire [31:0] s_0__15;
  wire [31:0] s_1__15;
  wire [1:0] S0__167;
  wire [10:0] S0__166;
  wire [8:0] S0__165;
  wire [9:0] S0__164;
  wire [31:0] and_58554;
  wire [31:0] S1__30;
  wire [31:0] value__43;
  wire [31:0] value__44;
  wire [31:0] S0__26;
  wire [31:0] maj__26;
  wire [31:0] temp1__121;
  wire [31:0] ch__30;
  wire [31:0] value__45;
  wire [31:0] temp2__26;
  wire [31:0] temp1__122;
  wire [31:0] temp1__288;
  wire [31:0] a__27;
  wire [31:0] temp1__124;
  wire [31:0] e__31;
  wire [2:0] s_0__111;
  wire [3:0] s_0__110;
  wire [10:0] s_0__109;
  wire [13:0] s_0__108;
  wire [9:0] s_1__111;
  wire [6:0] s_1__110;
  wire [1:0] s_1__109;
  wire [12:0] s_1__108;
  wire [5:0] S1__187;
  wire [4:0] S1__186;
  wire [13:0] S1__185;
  wire [6:0] S1__184;
  wire [31:0] s_0__16;
  wire [31:0] s_1__16;
  wire [1:0] S0__171;
  wire [10:0] S0__170;
  wire [8:0] S0__169;
  wire [9:0] S0__168;
  wire [31:0] and_58638;
  wire [31:0] S1__31;
  wire [31:0] value__46;
  wire [31:0] value__47;
  wire [31:0] S0__27;
  wire [31:0] maj__27;
  wire [31:0] temp1__125;
  wire [31:0] ch__31;
  wire [31:0] value__48;
  wire [31:0] temp2__27;
  wire [31:0] temp1__126;
  wire [31:0] temp1__289;
  wire [31:0] a__28;
  wire [31:0] temp1__128;
  wire [31:0] e__32;
  wire [2:0] s_0__115;
  wire [3:0] s_0__114;
  wire [10:0] s_0__113;
  wire [13:0] s_0__112;
  wire [9:0] s_1__115;
  wire [6:0] s_1__114;
  wire [1:0] s_1__113;
  wire [12:0] s_1__112;
  wire [5:0] S1__191;
  wire [4:0] S1__190;
  wire [13:0] S1__189;
  wire [6:0] S1__188;
  wire [31:0] s_0__17;
  wire [31:0] s_1__17;
  wire [1:0] S0__175;
  wire [10:0] S0__174;
  wire [8:0] S0__173;
  wire [9:0] S0__172;
  wire [31:0] and_58722;
  wire [31:0] S1__32;
  wire [31:0] value__49;
  wire [31:0] value__50;
  wire [31:0] S0__28;
  wire [31:0] maj__28;
  wire [31:0] temp1__129;
  wire [31:0] ch__32;
  wire [31:0] value__51;
  wire [2:0] s_0__119;
  wire [3:0] s_0__118;
  wire [10:0] s_0__117;
  wire [13:0] s_0__116;
  wire [9:0] s_1__119;
  wire [6:0] s_1__118;
  wire [1:0] s_1__117;
  wire [12:0] s_1__116;
  wire [31:0] temp2__28;
  wire [31:0] temp1__130;
  wire [31:0] temp1__290;
  wire [31:0] s_0__18;
  wire [31:0] s_1__18;
  wire [31:0] a__29;
  wire [31:0] temp1__132;
  wire [31:0] value__52;
  wire [31:0] value__53;
  wire [31:0] e__33;
  wire [31:0] value__54;
  wire [1:0] S0__179;
  wire [10:0] S0__178;
  wire [8:0] S0__177;
  wire [9:0] S0__176;
  wire [31:0] and_58807;
  wire [5:0] S1__195;
  wire [4:0] S1__194;
  wire [13:0] S1__193;
  wire [6:0] S1__192;
  wire [28:0] add_58815;
  wire [31:0] S0__29;
  wire [31:0] maj__29;
  wire [31:0] S1__33;
  wire [31:0] ch__33;
  wire [31:0] temp1__291;
  wire [2:0] s_0__123;
  wire [3:0] s_0__122;
  wire [10:0] s_0__121;
  wire [13:0] s_0__120;
  wire [9:0] s_1__123;
  wire [6:0] s_1__122;
  wire [1:0] s_1__121;
  wire [12:0] s_1__120;
  wire [31:0] temp2__29;
  wire [31:0] temp1__395;
  wire [31:0] temp1__396;
  wire [31:0] s_0__19;
  wire [31:0] s_1__19;
  wire [31:0] a__30;
  wire [31:0] temp1__397;
  wire [31:0] value__55;
  wire [31:0] value__56;
  wire [31:0] e__34;
  wire [31:0] value__57;
  wire [1:0] S0__183;
  wire [10:0] S0__182;
  wire [8:0] S0__181;
  wire [9:0] S0__180;
  wire [31:0] and_58894;
  wire [5:0] S1__199;
  wire [4:0] S1__198;
  wire [13:0] S1__197;
  wire [6:0] S1__196;
  wire [29:0] add_58902;
  wire [31:0] S0__30;
  wire [31:0] maj__30;
  wire [31:0] S1__34;
  wire [31:0] ch__34;
  wire [31:0] temp1__292;
  wire [31:0] temp2__30;
  wire [31:0] temp1__392;
  wire [31:0] temp1__393;
  wire [31:0] a__31;
  wire [31:0] temp1__394;
  wire [31:0] e__35;
  wire [2:0] s_0__127;
  wire [3:0] s_0__126;
  wire [10:0] s_0__125;
  wire [13:0] s_0__124;
  wire [9:0] s_1__127;
  wire [6:0] s_1__126;
  wire [1:0] s_1__125;
  wire [12:0] s_1__124;
  wire [5:0] S1__203;
  wire [4:0] S1__202;
  wire [13:0] S1__201;
  wire [6:0] S1__200;
  wire [31:0] s_0__20;
  wire [31:0] s_1__20;
  wire [1:0] S0__187;
  wire [10:0] S0__186;
  wire [8:0] S0__185;
  wire [9:0] S0__184;
  wire [31:0] and_58980;
  wire [31:0] S1__35;
  wire [31:0] value__58;
  wire [31:0] value__59;
  wire [31:0] S0__31;
  wire [31:0] maj__31;
  wire [31:0] temp1__141;
  wire [31:0] ch__35;
  wire [31:0] value__60;
  wire [2:0] s_0__131;
  wire [3:0] s_0__130;
  wire [10:0] s_0__129;
  wire [13:0] s_0__128;
  wire [9:0] s_1__131;
  wire [6:0] s_1__130;
  wire [1:0] s_1__129;
  wire [12:0] s_1__128;
  wire [31:0] temp2__31;
  wire [31:0] temp1__142;
  wire [31:0] temp1__293;
  wire [31:0] s_0__21;
  wire [31:0] s_1__21;
  wire [31:0] a__32;
  wire [31:0] temp1__144;
  wire [31:0] value__61;
  wire [31:0] value__62;
  wire [31:0] e__36;
  wire [31:0] value__63;
  wire [1:0] S0__191;
  wire [10:0] S0__190;
  wire [8:0] S0__189;
  wire [9:0] S0__188;
  wire [31:0] and_59064;
  wire [5:0] S1__207;
  wire [4:0] S1__206;
  wire [13:0] S1__205;
  wire [6:0] S1__204;
  wire [29:0] add_59072;
  wire [31:0] S0__32;
  wire [31:0] maj__32;
  wire [31:0] S1__36;
  wire [31:0] ch__36;
  wire [31:0] temp1__294;
  wire [31:0] temp2__32;
  wire [31:0] temp1__389;
  wire [31:0] temp1__390;
  wire [31:0] a__33;
  wire [31:0] temp1__391;
  wire [31:0] e__37;
  wire [2:0] s_0__135;
  wire [3:0] s_0__134;
  wire [10:0] s_0__133;
  wire [13:0] s_0__132;
  wire [9:0] s_1__135;
  wire [6:0] s_1__134;
  wire [1:0] s_1__133;
  wire [12:0] s_1__132;
  wire [5:0] S1__211;
  wire [4:0] S1__210;
  wire [13:0] S1__209;
  wire [6:0] S1__208;
  wire [31:0] s_0__22;
  wire [31:0] s_1__22;
  wire [1:0] S0__195;
  wire [10:0] S0__194;
  wire [8:0] S0__193;
  wire [9:0] S0__192;
  wire [31:0] and_59150;
  wire [31:0] S1__37;
  wire [31:0] value__64;
  wire [31:0] value__65;
  wire [31:0] S0__33;
  wire [31:0] maj__33;
  wire [31:0] temp1__149;
  wire [31:0] ch__37;
  wire [31:0] value__66;
  wire [2:0] s_0__139;
  wire [3:0] s_0__138;
  wire [10:0] s_0__137;
  wire [13:0] s_0__136;
  wire [9:0] s_1__139;
  wire [6:0] s_1__138;
  wire [1:0] s_1__137;
  wire [12:0] s_1__136;
  wire [31:0] temp2__33;
  wire [31:0] temp1__150;
  wire [31:0] temp1__295;
  wire [31:0] s_0__23;
  wire [31:0] s_1__23;
  wire [31:0] a__34;
  wire [31:0] temp1__152;
  wire [31:0] value__67;
  wire [31:0] value__68;
  wire [31:0] e__38;
  wire [31:0] value__69;
  wire [1:0] S0__199;
  wire [10:0] S0__198;
  wire [8:0] S0__197;
  wire [9:0] S0__196;
  wire [31:0] and_59234;
  wire [5:0] S1__215;
  wire [4:0] S1__214;
  wire [13:0] S1__213;
  wire [6:0] S1__212;
  wire [30:0] add_59242;
  wire [31:0] S0__34;
  wire [31:0] maj__34;
  wire [31:0] S1__38;
  wire [31:0] ch__38;
  wire [31:0] temp1__296;
  wire [31:0] temp2__34;
  wire [31:0] temp1__386;
  wire [31:0] temp1__387;
  wire [31:0] a__35;
  wire [31:0] temp1__388;
  wire [31:0] e__39;
  wire [2:0] s_0__143;
  wire [3:0] s_0__142;
  wire [10:0] s_0__141;
  wire [13:0] s_0__140;
  wire [9:0] s_1__143;
  wire [6:0] s_1__142;
  wire [1:0] s_1__141;
  wire [12:0] s_1__140;
  wire [5:0] S1__219;
  wire [4:0] S1__218;
  wire [13:0] S1__217;
  wire [6:0] S1__216;
  wire [31:0] s_0__24;
  wire [31:0] s_1__24;
  wire [1:0] S0__203;
  wire [10:0] S0__202;
  wire [8:0] S0__201;
  wire [9:0] S0__200;
  wire [31:0] and_59320;
  wire [31:0] S1__39;
  wire [31:0] value__70;
  wire [31:0] value__71;
  wire [31:0] S0__35;
  wire [31:0] maj__35;
  wire [31:0] temp1__157;
  wire [31:0] ch__39;
  wire [31:0] value__72;
  wire [31:0] temp2__35;
  wire [31:0] temp1__158;
  wire [31:0] temp1__297;
  wire [31:0] a__36;
  wire [31:0] temp1__160;
  wire [31:0] e__40;
  wire [2:0] s_0__147;
  wire [3:0] s_0__146;
  wire [10:0] s_0__145;
  wire [13:0] s_0__144;
  wire [9:0] s_1__147;
  wire [6:0] s_1__146;
  wire [1:0] s_1__145;
  wire [12:0] s_1__144;
  wire [5:0] S1__223;
  wire [4:0] S1__222;
  wire [13:0] S1__221;
  wire [6:0] S1__220;
  wire [31:0] s_0__25;
  wire [31:0] s_1__25;
  wire [1:0] S0__207;
  wire [10:0] S0__206;
  wire [8:0] S0__205;
  wire [9:0] S0__204;
  wire [31:0] and_59404;
  wire [31:0] S1__40;
  wire [31:0] value__73;
  wire [31:0] value__74;
  wire [31:0] S0__36;
  wire [31:0] maj__36;
  wire [31:0] temp1__161;
  wire [31:0] ch__40;
  wire [31:0] value__75;
  wire [31:0] temp2__36;
  wire [31:0] temp1__162;
  wire [31:0] temp1__298;
  wire [31:0] a__37;
  wire [31:0] temp1__164;
  wire [31:0] e__41;
  wire [2:0] s_0__151;
  wire [3:0] s_0__150;
  wire [10:0] s_0__149;
  wire [13:0] s_0__148;
  wire [9:0] s_1__151;
  wire [6:0] s_1__150;
  wire [1:0] s_1__149;
  wire [12:0] s_1__148;
  wire [5:0] S1__227;
  wire [4:0] S1__226;
  wire [13:0] S1__225;
  wire [6:0] S1__224;
  wire [31:0] s_0__26;
  wire [31:0] s_1__26;
  wire [1:0] S0__211;
  wire [10:0] S0__210;
  wire [8:0] S0__209;
  wire [9:0] S0__208;
  wire [31:0] and_59488;
  wire [31:0] S1__41;
  wire [31:0] value__76;
  wire [31:0] value__77;
  wire [31:0] S0__37;
  wire [31:0] maj__37;
  wire [31:0] temp1__165;
  wire [31:0] ch__41;
  wire [31:0] value__78;
  wire [2:0] s_0__155;
  wire [3:0] s_0__154;
  wire [10:0] s_0__153;
  wire [13:0] s_0__152;
  wire [9:0] s_1__155;
  wire [6:0] s_1__154;
  wire [1:0] s_1__153;
  wire [12:0] s_1__152;
  wire [31:0] temp2__37;
  wire [31:0] temp1__166;
  wire [31:0] temp1__299;
  wire [31:0] s_0__27;
  wire [31:0] s_1__27;
  wire [31:0] a__38;
  wire [31:0] temp1__168;
  wire [31:0] value__79;
  wire [31:0] value__80;
  wire [31:0] e__42;
  wire [31:0] value__81;
  wire [1:0] S0__215;
  wire [10:0] S0__214;
  wire [8:0] S0__213;
  wire [9:0] S0__212;
  wire [31:0] and_59573;
  wire [5:0] S1__231;
  wire [4:0] S1__230;
  wire [13:0] S1__229;
  wire [6:0] S1__228;
  wire [27:0] add_59581;
  wire [31:0] S0__38;
  wire [31:0] maj__38;
  wire [31:0] S1__42;
  wire [31:0] ch__42;
  wire [31:0] temp1__300;
  wire [31:0] temp2__38;
  wire [31:0] temp1__383;
  wire [31:0] temp1__384;
  wire [31:0] a__39;
  wire [31:0] temp1__385;
  wire [31:0] e__43;
  wire [2:0] s_0__159;
  wire [3:0] s_0__158;
  wire [10:0] s_0__157;
  wire [13:0] s_0__156;
  wire [9:0] s_1__159;
  wire [6:0] s_1__158;
  wire [1:0] s_1__157;
  wire [12:0] s_1__156;
  wire [5:0] S1__235;
  wire [4:0] S1__234;
  wire [13:0] S1__233;
  wire [6:0] S1__232;
  wire [31:0] s_0__28;
  wire [31:0] s_1__28;
  wire [1:0] S0__219;
  wire [10:0] S0__218;
  wire [8:0] S0__217;
  wire [9:0] S0__216;
  wire [31:0] and_59659;
  wire [31:0] S1__43;
  wire [31:0] value__82;
  wire [31:0] value__83;
  wire [31:0] S0__39;
  wire [31:0] maj__39;
  wire [31:0] temp1__173;
  wire [31:0] ch__43;
  wire [31:0] value__84;
  wire [31:0] temp2__39;
  wire [31:0] temp1__174;
  wire [31:0] temp1__301;
  wire [31:0] a__40;
  wire [31:0] temp1__176;
  wire [31:0] e__44;
  wire [2:0] s_0__163;
  wire [3:0] s_0__162;
  wire [10:0] s_0__161;
  wire [13:0] s_0__160;
  wire [9:0] s_1__163;
  wire [6:0] s_1__162;
  wire [1:0] s_1__161;
  wire [12:0] s_1__160;
  wire [5:0] S1__239;
  wire [4:0] S1__238;
  wire [13:0] S1__237;
  wire [6:0] S1__236;
  wire [31:0] s_0__29;
  wire [31:0] s_1__29;
  wire [1:0] S0__223;
  wire [10:0] S0__222;
  wire [8:0] S0__221;
  wire [9:0] S0__220;
  wire [31:0] and_59743;
  wire [31:0] S1__44;
  wire [31:0] value__85;
  wire [31:0] value__86;
  wire [31:0] S0__40;
  wire [31:0] maj__40;
  wire [31:0] temp1__177;
  wire [31:0] ch__44;
  wire [31:0] value__87;
  wire [2:0] s_0__167;
  wire [3:0] s_0__166;
  wire [10:0] s_0__165;
  wire [13:0] s_0__164;
  wire [9:0] s_1__167;
  wire [6:0] s_1__166;
  wire [1:0] s_1__165;
  wire [12:0] s_1__164;
  wire [31:0] temp2__40;
  wire [31:0] temp1__178;
  wire [31:0] temp1__302;
  wire [31:0] s_0__30;
  wire [31:0] s_1__30;
  wire [31:0] a__41;
  wire [31:0] temp1__180;
  wire [31:0] value__88;
  wire [31:0] value__89;
  wire [31:0] e__45;
  wire [31:0] value__90;
  wire [1:0] S0__227;
  wire [10:0] S0__226;
  wire [8:0] S0__225;
  wire [9:0] S0__224;
  wire [31:0] and_59828;
  wire [5:0] S1__243;
  wire [4:0] S1__242;
  wire [13:0] S1__241;
  wire [6:0] S1__240;
  wire [29:0] add_59836;
  wire [31:0] S0__41;
  wire [31:0] maj__41;
  wire [31:0] S1__45;
  wire [31:0] ch__45;
  wire [31:0] temp1__303;
  wire [31:0] temp2__41;
  wire [31:0] temp1__380;
  wire [31:0] temp1__381;
  wire [31:0] a__42;
  wire [31:0] temp1__382;
  wire [31:0] e__46;
  wire [2:0] s_0__171;
  wire [3:0] s_0__170;
  wire [10:0] s_0__169;
  wire [13:0] s_0__168;
  wire [9:0] s_1__171;
  wire [6:0] s_1__170;
  wire [1:0] s_1__169;
  wire [12:0] s_1__168;
  wire [5:0] S1__247;
  wire [4:0] S1__246;
  wire [13:0] S1__245;
  wire [6:0] S1__244;
  wire [31:0] s_0__31;
  wire [31:0] s_1__31;
  wire [1:0] S0__231;
  wire [10:0] S0__230;
  wire [8:0] S0__229;
  wire [9:0] S0__228;
  wire [31:0] and_59914;
  wire [31:0] S1__46;
  wire [31:0] value__91;
  wire [31:0] value__92;
  wire [31:0] S0__42;
  wire [31:0] maj__42;
  wire [31:0] temp1__185;
  wire [31:0] ch__46;
  wire [31:0] value__93;
  wire [2:0] s_0__175;
  wire [3:0] s_0__174;
  wire [10:0] s_0__173;
  wire [13:0] s_0__172;
  wire [9:0] s_1__175;
  wire [6:0] s_1__174;
  wire [1:0] s_1__173;
  wire [12:0] s_1__172;
  wire [31:0] temp2__42;
  wire [31:0] temp1__186;
  wire [31:0] temp1__304;
  wire [31:0] s_0__32;
  wire [31:0] s_1__32;
  wire [31:0] a__43;
  wire [31:0] temp1__188;
  wire [31:0] value__94;
  wire [31:0] value__95;
  wire [31:0] e__47;
  wire [31:0] value__96;
  wire [1:0] S0__235;
  wire [10:0] S0__234;
  wire [8:0] S0__233;
  wire [9:0] S0__232;
  wire [31:0] and_59998;
  wire [5:0] S1__251;
  wire [4:0] S1__250;
  wire [13:0] S1__249;
  wire [6:0] S1__248;
  wire [27:0] add_60006;
  wire [31:0] S0__43;
  wire [31:0] maj__43;
  wire [31:0] S1__47;
  wire [31:0] ch__47;
  wire [31:0] temp1__305;
  wire [2:0] s_0__179;
  wire [3:0] s_0__178;
  wire [10:0] s_0__177;
  wire [13:0] s_0__176;
  wire [9:0] s_1__179;
  wire [6:0] s_1__178;
  wire [1:0] s_1__177;
  wire [12:0] s_1__176;
  wire [31:0] temp2__43;
  wire [31:0] temp1__377;
  wire [31:0] temp1__378;
  wire [31:0] s_0__33;
  wire [31:0] s_1__33;
  wire [31:0] a__44;
  wire [31:0] temp1__379;
  wire [31:0] value__97;
  wire [31:0] value__98;
  wire [31:0] e__48;
  wire [31:0] value__99;
  wire [1:0] S0__239;
  wire [10:0] S0__238;
  wire [8:0] S0__237;
  wire [9:0] S0__236;
  wire [31:0] and_60085;
  wire [5:0] S1__255;
  wire [4:0] S1__254;
  wire [13:0] S1__253;
  wire [6:0] S1__252;
  wire [30:0] add_60093;
  wire [31:0] S0__44;
  wire [31:0] maj__44;
  wire [31:0] S1__48;
  wire [31:0] ch__48;
  wire [31:0] temp1__306;
  wire [2:0] s_0__183;
  wire [3:0] s_0__182;
  wire [10:0] s_0__181;
  wire [13:0] s_0__180;
  wire [9:0] s_1__183;
  wire [6:0] s_1__182;
  wire [1:0] s_1__181;
  wire [12:0] s_1__180;
  wire [31:0] temp2__44;
  wire [31:0] temp1__374;
  wire [31:0] temp1__375;
  wire [31:0] s_0__34;
  wire [31:0] s_1__34;
  wire [31:0] a__45;
  wire [31:0] temp1__376;
  wire [31:0] value__100;
  wire [31:0] value__101;
  wire [31:0] e__49;
  wire [31:0] value__102;
  wire [1:0] S0__243;
  wire [10:0] S0__242;
  wire [8:0] S0__241;
  wire [9:0] S0__240;
  wire [31:0] and_60172;
  wire [5:0] S1__259;
  wire [4:0] S1__258;
  wire [13:0] S1__257;
  wire [6:0] S1__256;
  wire [28:0] add_60180;
  wire [31:0] S0__45;
  wire [31:0] maj__45;
  wire [31:0] S1__49;
  wire [31:0] ch__49;
  wire [31:0] temp1__307;
  wire [2:0] s_0__187;
  wire [3:0] s_0__186;
  wire [10:0] s_0__185;
  wire [13:0] s_0__184;
  wire [9:0] s_1__187;
  wire [6:0] s_1__186;
  wire [1:0] s_1__185;
  wire [12:0] s_1__184;
  wire [31:0] temp2__45;
  wire [31:0] temp1__371;
  wire [31:0] temp1__372;
  wire [31:0] s_0__35;
  wire [31:0] s_1__35;
  wire [31:0] a__46;
  wire [31:0] temp1__373;
  wire [31:0] value__103;
  wire [31:0] value__104;
  wire [31:0] e__50;
  wire [31:0] value__105;
  wire [1:0] S0__247;
  wire [10:0] S0__246;
  wire [8:0] S0__245;
  wire [9:0] S0__244;
  wire [31:0] and_60259;
  wire [5:0] S1__263;
  wire [4:0] S1__262;
  wire [13:0] S1__261;
  wire [6:0] S1__260;
  wire [29:0] add_60267;
  wire [31:0] S0__46;
  wire [31:0] maj__46;
  wire [31:0] S1__50;
  wire [31:0] ch__50;
  wire [31:0] temp1__308;
  wire [31:0] temp2__46;
  wire [31:0] temp1__368;
  wire [31:0] temp1__369;
  wire [31:0] a__47;
  wire [31:0] temp1__370;
  wire [31:0] e__51;
  wire [2:0] s_0__191;
  wire [3:0] s_0__190;
  wire [10:0] s_0__189;
  wire [13:0] s_0__188;
  wire [9:0] s_1__191;
  wire [6:0] s_1__190;
  wire [1:0] s_1__189;
  wire [12:0] s_1__188;
  wire [5:0] S1__267;
  wire [4:0] S1__266;
  wire [13:0] S1__265;
  wire [6:0] S1__264;
  wire [31:0] s_0__36;
  wire [31:0] s_1__36;
  wire [1:0] S0__251;
  wire [10:0] S0__250;
  wire [8:0] S0__249;
  wire [9:0] S0__248;
  wire [31:0] and_60345;
  wire [31:0] S1__51;
  wire [31:0] value__106;
  wire [31:0] value__107;
  wire [31:0] S0__47;
  wire [31:0] maj__47;
  wire [31:0] temp1__205;
  wire [31:0] ch__51;
  wire [31:0] value__108;
  wire [31:0] temp2__47;
  wire [31:0] temp1__206;
  wire [31:0] temp1__309;
  wire [31:0] a__48;
  wire [31:0] temp1__208;
  wire [31:0] e__52;
  wire [2:0] s_0__195;
  wire [3:0] s_0__194;
  wire [10:0] s_0__193;
  wire [13:0] s_0__192;
  wire [9:0] s_1__195;
  wire [6:0] s_1__194;
  wire [1:0] s_1__193;
  wire [12:0] s_1__192;
  wire [5:0] S1__271;
  wire [4:0] S1__270;
  wire [13:0] S1__269;
  wire [6:0] S1__268;
  wire [31:0] s_0__37;
  wire [31:0] s_1__37;
  wire [1:0] S0__255;
  wire [10:0] S0__254;
  wire [8:0] S0__253;
  wire [9:0] S0__252;
  wire [31:0] and_60428;
  wire [31:0] S1__52;
  wire [31:0] value__109;
  wire [31:0] value__110;
  wire [31:0] S0__48;
  wire [31:0] maj__48;
  wire [31:0] temp1__209;
  wire [31:0] ch__52;
  wire [31:0] value__111;
  wire [2:0] s_0__199;
  wire [3:0] s_0__198;
  wire [10:0] s_0__197;
  wire [13:0] s_0__196;
  wire [9:0] s_1__199;
  wire [6:0] s_1__198;
  wire [1:0] s_1__197;
  wire [12:0] s_1__196;
  wire [31:0] temp2__48;
  wire [31:0] temp1__210;
  wire [31:0] temp1__310;
  wire [31:0] s_0__38;
  wire [31:0] s_1__38;
  wire [31:0] a__49;
  wire [31:0] temp1__212;
  wire [31:0] value__112;
  wire [31:0] value__113;
  wire [31:0] e__53;
  wire [31:0] value__114;
  wire [1:0] S0__259;
  wire [10:0] S0__258;
  wire [8:0] S0__257;
  wire [9:0] S0__256;
  wire [31:0] and_60498;
  wire [31:0] S0__49;
  wire [31:0] maj__49;
  wire [5:0] S1__275;
  wire [4:0] S1__274;
  wire [13:0] S1__273;
  wire [6:0] S1__272;
  wire [30:0] add_60523;
  wire [31:0] temp2__49;
  wire [31:0] S1__53;
  wire [31:0] ch__53;
  wire [31:0] temp1__311;
  wire [31:0] a__50;
  wire [31:0] temp1__365;
  wire [31:0] temp1__366;
  wire [31:0] temp1__367;
  wire [1:0] S0__263;
  wire [10:0] S0__262;
  wire [8:0] S0__261;
  wire [9:0] S0__260;
  wire [31:0] and_60549;
  wire [31:0] e__54;
  wire [31:0] S0__50;
  wire [31:0] maj__50;
  wire [2:0] s_0__203;
  wire [3:0] s_0__202;
  wire [10:0] s_0__201;
  wire [13:0] s_0__200;
  wire [9:0] s_1__203;
  wire [6:0] s_1__202;
  wire [1:0] s_1__201;
  wire [12:0] s_1__200;
  wire [31:0] temp2__50;
  wire [5:0] S1__279;
  wire [4:0] S1__278;
  wire [13:0] S1__277;
  wire [6:0] S1__276;
  wire [31:0] s_0__39;
  wire [31:0] s_1__39;
  wire [31:0] a__51;
  wire [31:0] S1__54;
  wire [31:0] value__115;
  wire [31:0] value__116;
  wire [31:0] temp1__217;
  wire [31:0] ch__54;
  wire [31:0] value__117;
  wire [1:0] S0__267;
  wire [10:0] S0__266;
  wire [8:0] S0__265;
  wire [9:0] S0__264;
  wire [31:0] and_60630;
  wire [31:0] temp1__218;
  wire [31:0] temp1__312;
  wire [31:0] S0__51;
  wire [31:0] maj__51;
  wire [31:0] temp1__220;
  wire [31:0] temp2__51;
  wire [31:0] e__55;
  wire [31:0] a__52;
  wire [2:0] s_0__207;
  wire [3:0] s_0__206;
  wire [10:0] s_0__205;
  wire [13:0] s_0__204;
  wire [9:0] s_1__207;
  wire [6:0] s_1__206;
  wire [1:0] s_1__205;
  wire [12:0] s_1__204;
  wire [5:0] S1__283;
  wire [4:0] S1__282;
  wire [13:0] S1__281;
  wire [6:0] S1__280;
  wire [31:0] s_0__40;
  wire [31:0] s_1__40;
  wire [1:0] S0__271;
  wire [10:0] S0__270;
  wire [8:0] S0__269;
  wire [9:0] S0__268;
  wire [31:0] and_60705;
  wire [31:0] S1__55;
  wire [31:0] value__118;
  wire [31:0] value__119;
  wire [31:0] S0__52;
  wire [31:0] maj__52;
  wire [31:0] temp1__221;
  wire [31:0] ch__55;
  wire [31:0] value__120;
  wire [2:0] s_0__211;
  wire [3:0] s_0__210;
  wire [10:0] s_0__209;
  wire [13:0] s_0__208;
  wire [9:0] s_1__211;
  wire [6:0] s_1__210;
  wire [1:0] s_1__209;
  wire [12:0] s_1__208;
  wire [31:0] temp2__52;
  wire [31:0] temp1__222;
  wire [31:0] temp1__313;
  wire [31:0] s_0__41;
  wire [31:0] s_1__41;
  wire [31:0] a__53;
  wire [31:0] temp1__224;
  wire [31:0] value__121;
  wire [31:0] value__122;
  wire [31:0] e__56;
  wire [31:0] value__123;
  wire [1:0] S0__275;
  wire [10:0] S0__274;
  wire [8:0] S0__273;
  wire [9:0] S0__272;
  wire [31:0] and_60775;
  wire [31:0] S0__53;
  wire [31:0] maj__53;
  wire [5:0] S1__287;
  wire [4:0] S1__286;
  wire [13:0] S1__285;
  wire [6:0] S1__284;
  wire [30:0] add_60800;
  wire [31:0] temp2__53;
  wire [31:0] S1__56;
  wire [31:0] ch__56;
  wire [31:0] temp1__314;
  wire [31:0] a__54;
  wire [31:0] temp1__362;
  wire [31:0] temp1__363;
  wire [31:0] temp1__364;
  wire [1:0] S0__279;
  wire [10:0] S0__278;
  wire [8:0] S0__277;
  wire [9:0] S0__276;
  wire [31:0] and_60826;
  wire [31:0] e__57;
  wire [31:0] S0__54;
  wire [31:0] maj__54;
  wire [2:0] s_0__215;
  wire [3:0] s_0__214;
  wire [10:0] s_0__213;
  wire [13:0] s_0__212;
  wire [9:0] s_1__215;
  wire [6:0] s_1__214;
  wire [1:0] s_1__213;
  wire [12:0] s_1__212;
  wire [31:0] temp2__54;
  wire [5:0] S1__291;
  wire [4:0] S1__290;
  wire [13:0] S1__289;
  wire [6:0] S1__288;
  wire [31:0] s_0__42;
  wire [31:0] s_1__42;
  wire [31:0] a__55;
  wire [31:0] S1__57;
  wire [31:0] value__124;
  wire [31:0] value__125;
  wire [31:0] temp1__229;
  wire [31:0] ch__57;
  wire [31:0] value__126;
  wire [2:0] s_0__219;
  wire [3:0] s_0__218;
  wire [10:0] s_0__217;
  wire [13:0] s_0__216;
  wire [9:0] s_1__219;
  wire [6:0] s_1__218;
  wire [1:0] s_1__217;
  wire [12:0] s_1__216;
  wire [1:0] S0__283;
  wire [10:0] S0__282;
  wire [8:0] S0__281;
  wire [9:0] S0__280;
  wire [31:0] and_60936;
  wire [31:0] temp1__230;
  wire [31:0] temp1__315;
  wire [31:0] s_0__43;
  wire [31:0] s_1__43;
  wire [31:0] S0__55;
  wire [31:0] maj__55;
  wire [31:0] temp1__232;
  wire [31:0] value__127;
  wire [31:0] value__128;
  wire [31:0] temp2__55;
  wire [31:0] e__58;
  wire [31:0] value__129;
  wire [31:0] a__56;
  wire [5:0] S1__295;
  wire [4:0] S1__294;
  wire [13:0] S1__293;
  wire [6:0] S1__292;
  wire [29:0] add_60984;
  wire [1:0] S0__287;
  wire [10:0] S0__286;
  wire [8:0] S0__285;
  wire [9:0] S0__284;
  wire [31:0] and_61012;
  wire [31:0] S1__58;
  wire [31:0] ch__58;
  wire [31:0] temp1__316;
  wire [2:0] s_0__223;
  wire [3:0] s_0__222;
  wire [10:0] s_0__221;
  wire [13:0] s_0__220;
  wire [9:0] s_1__223;
  wire [6:0] s_1__222;
  wire [1:0] s_1__221;
  wire [12:0] s_1__220;
  wire [31:0] S0__56;
  wire [31:0] maj__56;
  wire [31:0] temp1__359;
  wire [31:0] temp1__360;
  wire [31:0] s_0__44;
  wire [31:0] s_1__44;
  wire [31:0] temp2__56;
  wire [31:0] temp1__361;
  wire [31:0] value__130;
  wire [31:0] value__131;
  wire [31:0] a__57;
  wire [31:0] e__59;
  wire [31:0] value__132;
  wire [1:0] S0__291;
  wire [10:0] S0__290;
  wire [8:0] S0__289;
  wire [9:0] S0__288;
  wire [31:0] and_61069;
  wire [5:0] S1__299;
  wire [4:0] S1__298;
  wire [13:0] S1__297;
  wire [6:0] S1__296;
  wire [28:0] add_61077;
  wire [31:0] S0__57;
  wire [31:0] maj__57;
  wire [31:0] S1__59;
  wire [31:0] ch__59;
  wire [31:0] temp1__317;
  wire [2:0] s_0__227;
  wire [3:0] s_0__226;
  wire [10:0] s_0__225;
  wire [13:0] s_0__224;
  wire [9:0] s_1__227;
  wire [6:0] s_1__226;
  wire [1:0] s_1__225;
  wire [12:0] s_1__224;
  wire [31:0] temp2__57;
  wire [31:0] temp1__356;
  wire [31:0] temp1__357;
  wire [31:0] s_0__45;
  wire [31:0] s_1__45;
  wire [31:0] a__58;
  wire [31:0] temp1__358;
  wire [31:0] value__133;
  wire [31:0] value__134;
  wire [31:0] e__60;
  wire [31:0] value__135;
  wire [1:0] S0__295;
  wire [10:0] S0__294;
  wire [8:0] S0__293;
  wire [9:0] S0__292;
  wire [31:0] and_61140;
  wire [31:0] S0__58;
  wire [31:0] maj__58;
  wire [5:0] S1__303;
  wire [4:0] S1__302;
  wire [13:0] S1__301;
  wire [6:0] S1__300;
  wire [30:0] add_61165;
  wire [31:0] temp2__58;
  wire [31:0] S1__60;
  wire [31:0] ch__60;
  wire [31:0] temp1__318;
  wire [31:0] a__59;
  wire [31:0] temp1__353;
  wire [31:0] temp1__354;
  wire [31:0] temp1__355;
  wire [1:0] S0__299;
  wire [10:0] S0__298;
  wire [8:0] S0__297;
  wire [9:0] S0__296;
  wire [31:0] and_61191;
  wire [31:0] e__61;
  wire [31:0] S0__59;
  wire [31:0] maj__59;
  wire [2:0] s_0__231;
  wire [3:0] s_0__230;
  wire [10:0] s_0__229;
  wire [13:0] s_0__228;
  wire [9:0] s_1__231;
  wire [6:0] s_1__230;
  wire [1:0] s_1__229;
  wire [12:0] s_1__228;
  wire [31:0] temp2__59;
  wire [5:0] S1__307;
  wire [4:0] S1__306;
  wire [13:0] S1__305;
  wire [6:0] S1__304;
  wire [31:0] s_0__46;
  wire [31:0] s_1__46;
  wire [31:0] a__60;
  wire [31:0] S1__61;
  wire [31:0] value__136;
  wire [31:0] value__137;
  wire [31:0] temp1__245;
  wire [31:0] ch__61;
  wire [31:0] value__138;
  wire [1:0] S0__303;
  wire [10:0] S0__302;
  wire [8:0] S0__301;
  wire [9:0] S0__300;
  wire [31:0] and_61272;
  wire [31:0] temp1__246;
  wire [31:0] temp1__319;
  wire [31:0] S0__60;
  wire [31:0] maj__60;
  wire [31:0] temp1__248;
  wire [31:0] temp2__60;
  wire [31:0] e__62;
  wire [31:0] a__61;
  wire [5:0] S1__311;
  wire [4:0] S1__310;
  wire [13:0] S1__309;
  wire [6:0] S1__308;
  wire [2:0] s_0__235;
  wire [3:0] s_0__234;
  wire [10:0] s_0__233;
  wire [13:0] s_0__232;
  wire [9:0] s_1__235;
  wire [6:0] s_1__234;
  wire [1:0] s_1__233;
  wire [12:0] s_1__232;
  wire [1:0] S0__307;
  wire [10:0] S0__306;
  wire [8:0] S0__305;
  wire [9:0] S0__304;
  wire [31:0] and_61346;
  wire [31:0] S1__62;
  wire [31:0] ch__62;
  wire [31:0] s_0__47;
  wire [31:0] s_1__47;
  wire [31:0] S0__61;
  wire [31:0] maj__61;
  wire [31:0] temp1__346;
  wire [31:0] temp1__347;
  wire [31:0] temp1__348;
  wire [31:0] temp1__349;
  wire [31:0] temp2__61;
  wire [31:0] temp1__350;
  wire [31:0] temp1__351;
  wire [31:0] a__62;
  wire [31:0] temp1__352;
  wire [31:0] e__63;
  wire [12:0] s_1__236;
  wire [1:0] S0__311;
  wire [10:0] S0__310;
  wire [8:0] S0__309;
  wire [9:0] S0__308;
  wire [31:0] and_61393;
  wire [9:0] s_1__239;
  wire [6:0] s_1__238;
  wire [1:0] s_1__237;
  wire [31:0] S0__62;
  wire [31:0] maj__62;
  wire [5:0] S1__315;
  wire [4:0] S1__314;
  wire [13:0] S1__313;
  wire [6:0] S1__312;
  wire [2:0] s_0__239;
  wire [3:0] s_0__238;
  wire [10:0] s_0__237;
  wire [13:0] s_0__236;
  wire [31:0] temp2__62;
  wire [31:0] S1__63;
  wire [31:0] ch__63;
  wire [31:0] s_0__240;
  wire [30:0] add_61441;
  wire [31:0] a__63;
  wire [31:0] temp1__339;
  wire [31:0] temp1__340;
  wire [31:0] temp1__341;
  wire [31:0] temp1__342;
  wire [31:0] temp1__343;
  wire [31:0] temp1__344;
  wire [1:0] S0__315;
  wire [10:0] S0__314;
  wire [8:0] S0__313;
  wire [9:0] S0__312;
  wire [31:0] temp1__345;
  wire [31:0] S0__63;
  wire [31:0] maj__63;
  wire [31:0] b__68;
  wire [31:0] add_61478;
  wire [31:0] add_61479;
  wire [31:0] c__66;
  wire [30:0] add_61481;
  wire [30:0] add_61483;
  wire [31:0] e__64;
  wire [31:0] f__66;
  wire [29:0] add_61487;
  wire [31:0] h__1;
  wire [31:0] h7;
  wire [31:0] add_61491;
  wire [31:0] add_61492;
  wire [31:0] add_61495;
  wire [31:0] add_61497;
  wire [31:0] add_61498;
  assign add_56574 = message[511:483] + 29'h1e6e_fdad;
  assign add_56578 = {add_56574, message[482:481]} + 31'h52a7_fa9d;
  assign e__66 = {add_56578, message[480]};
  assign f__1 = 32'h510e_527f;
  assign S1__67 = {add_56578[4:0], message[480]} ^ add_56578[9:4] ^ add_56578[23:18];
  assign S1__66 = add_56578[30:26] ^ {add_56578[3:0], message[480]} ^ add_56578[17:13];
  assign S1__65 = add_56578[25:12] ^ add_56578[30:17] ^ {add_56578[12:0], message[480]};
  assign S1__64 = add_56578[11:5] ^ add_56578[16:10] ^ add_56578[30:24];
  assign S1__1 = {S1__67, S1__66, S1__65, S1__64};
  assign ch__1 = e__66 & f__1 ^ ~(e__66 | 32'h64fa_9773);
  assign add_56608 = message[479:450] + 30'h242e_c78f;
  assign temp1__336 = S1__1 + ch__1;
  assign temp1__337 = {add_56608, message[449:448]};
  assign temp1__338 = temp1__336 + temp1__337;
  assign add_56615 = temp1__338[31:1] + 31'h1e37_79b9;
  assign e__67 = {add_56615, temp1__338[0]};
  assign S1__71 = {add_56615[4:0], temp1__338[0]} ^ add_56615[9:4] ^ add_56615[23:18];
  assign S1__70 = add_56615[30:26] ^ {add_56615[3:0], temp1__338[0]} ^ add_56615[17:13];
  assign S1__69 = add_56615[25:12] ^ add_56615[30:17] ^ {add_56615[12:0], temp1__338[0]};
  assign S1__68 = add_56615[11:5] ^ add_56615[16:10] ^ add_56615[30:24];
  assign S1__2 = {S1__71, S1__70, S1__69, S1__68};
  assign ch__2 = {add_56615 & add_56578, temp1__338[0] & message[480]} ^ ~(e__67 | 32'haef1_ad80);
  assign w_im15__1 = message[447:416];
  assign temp1__331 = 32'h50c6_645b;
  assign temp1__332 = S1__2 + ch__2;
  assign temp1__333 = w_im15__1 + temp1__331;
  assign temp1__334 = temp1__332 + temp1__333;
  assign c__67 = 32'hbb67_ae85;
  assign e__68 = temp1__334 + c__67;
  assign S1__75 = e__68[5:0] ^ e__68[10:5] ^ e__68[24:19];
  assign S1__74 = e__68[31:27] ^ e__68[4:0] ^ e__68[18:14];
  assign S1__73 = e__68[26:13] ^ e__68[31:18] ^ e__68[13:0];
  assign S1__72 = e__68[12:6] ^ e__68[17:11] ^ e__68[31:25];
  assign S1__3 = {S1__75, S1__74, S1__73, S1__72};
  assign ch__3 = e__68 & e__67 ^ ~(e__68 | {~add_56578, ~message[480]});
  assign add_56676 = message[415:386] + 30'h0eb1_0b89;
  assign temp1__328 = S1__3 + ch__3;
  assign temp1__329 = {add_56676, message[385:384]};
  assign temp1__330 = temp1__328 + temp1__329;
  assign b__67 = 32'h6a09_e667;
  assign e__69 = temp1__330 + b__67;
  assign S1__79 = e__69[5:0] ^ e__69[10:5] ^ e__69[24:19];
  assign S1__78 = e__69[31:27] ^ e__69[4:0] ^ e__69[18:14];
  assign S1__77 = e__69[26:13] ^ e__69[31:18] ^ e__69[13:0];
  assign S1__76 = e__69[12:6] ^ e__69[17:11] ^ e__69[31:25];
  assign S1__4 = {S1__79, S1__78, S1__77, S1__76};
  assign temp1__17 = e__66 + S1__4;
  assign ch__4 = e__69 & e__68 ^ ~(e__69 | {~add_56615, ~temp1__338[0]});
  assign w_im15__3 = message[383:352];
  assign temp1__323 = {add_56574, message[482:480]};
  assign temp2 = 32'h0890_9ae5;
  assign temp1__18 = temp1__17 + ch__4;
  assign temp1__262 = w_im15__3 + 32'h3956_c25b;
  assign a__1 = temp1__323 + temp2;
  assign temp1__20 = temp1__18 + temp1__262;
  assign e__5 = a__1 + temp1__20;
  assign b__1 = 32'h6a09_e667;
  assign c__1 = 32'hbb67_ae85;
  assign S1__83 = e__5[5:0] ^ e__5[10:5] ^ e__5[24:19];
  assign S1__82 = e__5[31:27] ^ e__5[4:0] ^ e__5[18:14];
  assign S1__81 = e__5[26:13] ^ e__5[31:18] ^ e__5[13:0];
  assign S1__80 = e__5[12:6] ^ e__5[17:11] ^ e__5[31:25];
  assign S0__67 = a__1[1:0] ^ a__1[12:11] ^ a__1[21:20];
  assign S0__66 = a__1[31:21] ^ a__1[10:0] ^ a__1[19:9];
  assign S0__65 = a__1[20:12] ^ a__1[31:23] ^ a__1[8:0];
  assign S0__64 = a__1[11:2] ^ a__1[22:13] ^ a__1[31:22];
  assign and_56752 = a__1 & b__1;
  assign S1__5 = {S1__83, S1__82, S1__81, S1__80};
  assign S0__1 = {S0__67, S0__66, S0__65, S0__64};
  assign maj__1 = and_56752 ^ a__1 & c__1 ^ 32'h2a01_a605;
  assign temp1__21 = e__67 + S1__5;
  assign ch__5 = e__5 & e__69 ^ ~(e__5 | ~e__68);
  assign w_im15__4 = message[351:320];
  assign temp2__1 = S0__1 + maj__1;
  assign temp1__22 = temp1__21 + ch__5;
  assign temp1__263 = w_im15__4 + 32'h59f1_11f1;
  assign a__2 = temp1__338 + temp2__1;
  assign temp1__24 = temp1__22 + temp1__263;
  assign e__6 = a__2 + temp1__24;
  assign b__66 = 32'h6a09_e667;
  assign S0__71 = a__2[1:0] ^ a__2[12:11] ^ a__2[21:20];
  assign S0__70 = a__2[31:21] ^ a__2[10:0] ^ a__2[19:9];
  assign S0__69 = a__2[20:12] ^ a__2[31:23] ^ a__2[8:0];
  assign S0__68 = a__2[11:2] ^ a__2[22:13] ^ a__2[31:22];
  assign and_56802 = a__2 & a__1;
  assign S1__87 = e__6[5:0] ^ e__6[10:5] ^ e__6[24:19];
  assign S1__86 = e__6[31:27] ^ e__6[4:0] ^ e__6[18:14];
  assign S1__85 = e__6[26:13] ^ e__6[31:18] ^ e__6[13:0];
  assign S1__84 = e__6[12:6] ^ e__6[17:11] ^ e__6[31:25];
  assign add_56810 = message[319:290] + 30'h248f_e0a9;
  assign S0__2 = {S0__71, S0__70, S0__69, S0__68};
  assign maj__2 = and_56802 ^ a__2 & b__66 ^ and_56752;
  assign S1__6 = {S1__87, S1__86, S1__85, S1__84};
  assign ch__6 = e__6 & e__5 ^ ~(e__6 | ~e__69);
  assign temp1__264 = {add_56810, message[289:288]};
  assign temp2__2 = S0__2 + maj__2;
  assign temp1__437 = e__68 + S1__6;
  assign temp1__438 = ch__6 + temp1__264;
  assign a__3 = temp1__334 + temp2__2;
  assign temp1__439 = temp1__437 + temp1__438;
  assign e__7 = a__3 + temp1__439;
  assign S1__91 = e__7[5:0] ^ e__7[10:5] ^ e__7[24:19];
  assign S1__90 = e__7[31:27] ^ e__7[4:0] ^ e__7[18:14];
  assign S1__89 = e__7[26:13] ^ e__7[31:18] ^ e__7[13:0];
  assign S1__88 = e__7[12:6] ^ e__7[17:11] ^ e__7[31:25];
  assign S0__75 = a__3[1:0] ^ a__3[12:11] ^ a__3[21:20];
  assign S0__74 = a__3[31:21] ^ a__3[10:0] ^ a__3[19:9];
  assign S0__73 = a__3[20:12] ^ a__3[31:23] ^ a__3[8:0];
  assign S0__72 = a__3[11:2] ^ a__3[22:13] ^ a__3[31:22];
  assign and_56856 = a__3 & a__2;
  assign S1__7 = {S1__91, S1__90, S1__89, S1__88};
  assign S0__3 = {S0__75, S0__74, S0__73, S0__72};
  assign maj__3 = and_56856 ^ a__3 & a__1 ^ and_56802;
  assign temp1__29 = e__69 + S1__7;
  assign ch__7 = e__7 & e__6 ^ ~(e__7 | ~e__5);
  assign w_im15__6 = message[287:256];
  assign temp2__3 = S0__3 + maj__3;
  assign temp1__30 = temp1__29 + ch__7;
  assign temp1__265 = w_im15__6 + 32'hab1c_5ed5;
  assign a__4 = temp1__330 + temp2__3;
  assign temp1__32 = temp1__30 + temp1__265;
  assign e__8 = a__4 + temp1__32;
  assign S0__79 = a__4[1:0] ^ a__4[12:11] ^ a__4[21:20];
  assign S0__78 = a__4[31:21] ^ a__4[10:0] ^ a__4[19:9];
  assign S0__77 = a__4[20:12] ^ a__4[31:23] ^ a__4[8:0];
  assign S0__76 = a__4[11:2] ^ a__4[22:13] ^ a__4[31:22];
  assign and_56904 = a__4 & a__3;
  assign S1__95 = e__8[5:0] ^ e__8[10:5] ^ e__8[24:19];
  assign S1__94 = e__8[31:27] ^ e__8[4:0] ^ e__8[18:14];
  assign S1__93 = e__8[26:13] ^ e__8[31:18] ^ e__8[13:0];
  assign S1__92 = e__8[12:6] ^ e__8[17:11] ^ e__8[31:25];
  assign add_56912 = message[255:227] + 29'h1b00_f553;
  assign S0__4 = {S0__79, S0__78, S0__77, S0__76};
  assign maj__4 = and_56904 ^ a__4 & a__2 ^ and_56856;
  assign S1__8 = {S1__95, S1__94, S1__93, S1__92};
  assign ch__8 = e__8 & e__7 ^ ~(e__8 | ~e__6);
  assign temp1__266 = {add_56912, message[226:224]};
  assign temp2__4 = S0__4 + maj__4;
  assign temp1__434 = e__5 + S1__8;
  assign temp1__435 = ch__8 + temp1__266;
  assign a__5 = temp1__20 + temp2__4;
  assign temp1__436 = temp1__434 + temp1__435;
  assign e__9 = a__5 + temp1__436;
  assign S1__99 = e__9[5:0] ^ e__9[10:5] ^ e__9[24:19];
  assign S1__98 = e__9[31:27] ^ e__9[4:0] ^ e__9[18:14];
  assign S1__97 = e__9[26:13] ^ e__9[31:18] ^ e__9[13:0];
  assign S1__96 = e__9[12:6] ^ e__9[17:11] ^ e__9[31:25];
  assign S0__83 = a__5[1:0] ^ a__5[12:11] ^ a__5[21:20];
  assign S0__82 = a__5[31:21] ^ a__5[10:0] ^ a__5[19:9];
  assign S0__81 = a__5[20:12] ^ a__5[31:23] ^ a__5[8:0];
  assign S0__80 = a__5[11:2] ^ a__5[22:13] ^ a__5[31:22];
  assign and_56958 = a__5 & a__4;
  assign S1__9 = {S1__99, S1__98, S1__97, S1__96};
  assign S0__5 = {S0__83, S0__82, S0__81, S0__80};
  assign maj__5 = and_56958 ^ a__5 & a__3 ^ and_56904;
  assign temp1__37 = e__6 + S1__9;
  assign ch__9 = e__9 & e__8 ^ ~(e__9 | ~e__7);
  assign w_im15__8 = message[223:192];
  assign temp2__5 = S0__5 + maj__5;
  assign temp1__38 = temp1__37 + ch__9;
  assign temp1__267 = w_im15__8 + 32'h1283_5b01;
  assign a__6 = temp1__24 + temp2__5;
  assign temp1__40 = temp1__38 + temp1__267;
  assign e__10 = a__6 + temp1__40;
  assign S0__87 = a__6[1:0] ^ a__6[12:11] ^ a__6[21:20];
  assign S0__86 = a__6[31:21] ^ a__6[10:0] ^ a__6[19:9];
  assign S0__85 = a__6[20:12] ^ a__6[31:23] ^ a__6[8:0];
  assign S0__84 = a__6[11:2] ^ a__6[22:13] ^ a__6[31:22];
  assign and_57006 = a__6 & a__5;
  assign S1__103 = e__10[5:0] ^ e__10[10:5] ^ e__10[24:19];
  assign S1__102 = e__10[31:27] ^ e__10[4:0] ^ e__10[18:14];
  assign S1__101 = e__10[26:13] ^ e__10[31:18] ^ e__10[13:0];
  assign S1__100 = e__10[12:6] ^ e__10[17:11] ^ e__10[31:25];
  assign add_57014 = message[191:161] + 31'h1218_c2df;
  assign S0__6 = {S0__87, S0__86, S0__85, S0__84};
  assign maj__6 = and_57006 ^ a__6 & a__4 ^ and_56958;
  assign S1__10 = {S1__103, S1__102, S1__101, S1__100};
  assign ch__10 = e__10 & e__9 ^ ~(e__10 | ~e__8);
  assign temp1__268 = {add_57014, message[160]};
  assign temp2__6 = S0__6 + maj__6;
  assign temp1__431 = e__7 + S1__10;
  assign temp1__432 = ch__10 + temp1__268;
  assign a__7 = temp1__439 + temp2__6;
  assign temp1__433 = temp1__431 + temp1__432;
  assign e__11 = a__7 + temp1__433;
  assign S1__107 = e__11[5:0] ^ e__11[10:5] ^ e__11[24:19];
  assign S1__106 = e__11[31:27] ^ e__11[4:0] ^ e__11[18:14];
  assign S1__105 = e__11[26:13] ^ e__11[31:18] ^ e__11[13:0];
  assign S1__104 = e__11[12:6] ^ e__11[17:11] ^ e__11[31:25];
  assign S0__91 = a__7[1:0] ^ a__7[12:11] ^ a__7[21:20];
  assign S0__90 = a__7[31:21] ^ a__7[10:0] ^ a__7[19:9];
  assign S0__89 = a__7[20:12] ^ a__7[31:23] ^ a__7[8:0];
  assign S0__88 = a__7[11:2] ^ a__7[22:13] ^ a__7[31:22];
  assign and_57060 = a__7 & a__6;
  assign S1__11 = {S1__107, S1__106, S1__105, S1__104};
  assign S0__7 = {S0__91, S0__90, S0__89, S0__88};
  assign maj__7 = and_57060 ^ a__7 & a__5 ^ and_57006;
  assign temp1__45 = e__8 + S1__11;
  assign ch__11 = e__11 & e__10 ^ ~(e__11 | ~e__9);
  assign w_im15__10 = message[159:128];
  assign temp2__7 = S0__7 + maj__7;
  assign temp1__46 = temp1__45 + ch__11;
  assign temp1__269 = w_im15__10 + 32'h550c_7dc3;
  assign a__8 = temp1__32 + temp2__7;
  assign temp1__48 = temp1__46 + temp1__269;
  assign e__12 = a__8 + temp1__48;
  assign S0__95 = a__8[1:0] ^ a__8[12:11] ^ a__8[21:20];
  assign S0__94 = a__8[31:21] ^ a__8[10:0] ^ a__8[19:9];
  assign S0__93 = a__8[20:12] ^ a__8[31:23] ^ a__8[8:0];
  assign S0__92 = a__8[11:2] ^ a__8[22:13] ^ a__8[31:22];
  assign and_57108 = a__8 & a__7;
  assign S1__111 = e__12[5:0] ^ e__12[10:5] ^ e__12[24:19];
  assign S1__110 = e__12[31:27] ^ e__12[4:0] ^ e__12[18:14];
  assign S1__109 = e__12[26:13] ^ e__12[31:18] ^ e__12[13:0];
  assign S1__108 = e__12[12:6] ^ e__12[17:11] ^ e__12[31:25];
  assign add_57116 = message[127:98] + 30'h1caf_975d;
  assign S0__8 = {S0__95, S0__94, S0__93, S0__92};
  assign maj__8 = and_57108 ^ a__8 & a__6 ^ and_57060;
  assign S1__12 = {S1__111, S1__110, S1__109, S1__108};
  assign ch__12 = e__12 & e__11 ^ ~(e__12 | ~e__10);
  assign temp1__270 = {add_57116, message[97:96]};
  assign temp2__8 = S0__8 + maj__8;
  assign temp1__428 = e__9 + S1__12;
  assign temp1__429 = ch__12 + temp1__270;
  assign a__9 = temp1__436 + temp2__8;
  assign temp1__430 = temp1__428 + temp1__429;
  assign e__13 = a__9 + temp1__430;
  assign S0__99 = a__9[1:0] ^ a__9[12:11] ^ a__9[21:20];
  assign S0__98 = a__9[31:21] ^ a__9[10:0] ^ a__9[19:9];
  assign S0__97 = a__9[20:12] ^ a__9[31:23] ^ a__9[8:0];
  assign S0__96 = a__9[11:2] ^ a__9[22:13] ^ a__9[31:22];
  assign and_57160 = a__9 & a__8;
  assign S1__115 = e__13[5:0] ^ e__13[10:5] ^ e__13[24:19];
  assign S1__114 = e__13[31:27] ^ e__13[4:0] ^ e__13[18:14];
  assign S1__113 = e__13[26:13] ^ e__13[31:18] ^ e__13[13:0];
  assign S1__112 = e__13[12:6] ^ e__13[17:11] ^ e__13[31:25];
  assign add_57168 = message[95:65] + 31'h406f_58ff;
  assign S0__9 = {S0__99, S0__98, S0__97, S0__96};
  assign maj__9 = and_57160 ^ a__9 & a__7 ^ and_57108;
  assign S1__13 = {S1__115, S1__114, S1__113, S1__112};
  assign ch__13 = e__13 & e__12 ^ ~(e__13 | ~e__11);
  assign temp1__271 = {add_57168, message[64]};
  assign temp2__9 = S0__9 + maj__9;
  assign temp1__425 = e__10 + S1__13;
  assign temp1__426 = ch__13 + temp1__271;
  assign a__10 = temp1__40 + temp2__9;
  assign temp1__427 = temp1__425 + temp1__426;
  assign e__14 = a__10 + temp1__427;
  assign S1__119 = e__14[5:0] ^ e__14[10:5] ^ e__14[24:19];
  assign S1__118 = e__14[31:27] ^ e__14[4:0] ^ e__14[18:14];
  assign S1__117 = e__14[26:13] ^ e__14[31:18] ^ e__14[13:0];
  assign S1__116 = e__14[12:6] ^ e__14[17:11] ^ e__14[31:25];
  assign S0__103 = a__10[1:0] ^ a__10[12:11] ^ a__10[21:20];
  assign S0__102 = a__10[31:21] ^ a__10[10:0] ^ a__10[19:9];
  assign S0__101 = a__10[20:12] ^ a__10[31:23] ^ a__10[8:0];
  assign S0__100 = a__10[11:2] ^ a__10[22:13] ^ a__10[31:22];
  assign and_57214 = a__10 & a__9;
  assign S1__14 = {S1__119, S1__118, S1__117, S1__116};
  assign S0__10 = {S0__103, S0__102, S0__101, S0__100};
  assign maj__10 = and_57214 ^ a__10 & a__8 ^ and_57160;
  assign temp1__57 = e__11 + S1__14;
  assign ch__14 = e__14 & e__13 ^ ~(e__14 | ~e__12);
  assign w_init_im2 = message[63:32];
  assign temp2__10 = S0__10 + maj__10;
  assign temp1__58 = temp1__57 + ch__14;
  assign temp1__272 = w_init_im2 + 32'h9bdc_06a7;
  assign a__11 = temp1__433 + temp2__10;
  assign temp1__60 = temp1__58 + temp1__272;
  assign e__15 = a__11 + temp1__60;
  assign S0__107 = a__11[1:0] ^ a__11[12:11] ^ a__11[21:20];
  assign S0__106 = a__11[31:21] ^ a__11[10:0] ^ a__11[19:9];
  assign S0__105 = a__11[20:12] ^ a__11[31:23] ^ a__11[8:0];
  assign S0__104 = a__11[11:2] ^ a__11[22:13] ^ a__11[31:22];
  assign and_57262 = a__11 & a__10;
  assign S1__123 = e__15[5:0] ^ e__15[10:5] ^ e__15[24:19];
  assign S1__122 = e__15[31:27] ^ e__15[4:0] ^ e__15[18:14];
  assign S1__121 = e__15[26:13] ^ e__15[31:18] ^ e__15[13:0];
  assign S1__120 = e__15[12:6] ^ e__15[17:11] ^ e__15[31:25];
  assign add_57270 = message[31:2] + 30'h3066_fc5d;
  assign S0__11 = {S0__107, S0__106, S0__105, S0__104};
  assign maj__11 = and_57262 ^ a__11 & a__9 ^ and_57214;
  assign S1__15 = {S1__123, S1__122, S1__121, S1__120};
  assign ch__15 = e__15 & e__14 ^ ~(e__15 | ~e__13);
  assign temp1__273 = {add_57270, message[1:0]};
  assign temp2__11 = S0__11 + maj__11;
  assign temp1__422 = e__12 + S1__15;
  assign temp1__423 = ch__15 + temp1__273;
  assign a__12 = temp1__48 + temp2__11;
  assign temp1__424 = temp1__422 + temp1__423;
  assign e__16 = a__12 + temp1__424;
  assign s_0__51 = message[454:452] ^ message[465:463];
  assign s_0__50 = message[451:448] ^ message[462:459] ^ message[479:476];
  assign s_0__49 = message[479:469] ^ message[458:448] ^ message[475:465];
  assign s_0__48 = message[468:455] ^ message[479:466] ^ message[464:451];
  assign s_1__51 = message[48:39] ^ message[50:41];
  assign s_1__50 = message[38:32] ^ message[40:34] ^ message[63:57];
  assign s_1__49 = message[63:62] ^ message[33:32] ^ message[56:55];
  assign s_1__48 = message[61:49] ^ message[63:51] ^ message[54:42];
  assign S1__127 = e__16[5:0] ^ e__16[10:5] ^ e__16[24:19];
  assign S1__126 = e__16[31:27] ^ e__16[4:0] ^ e__16[18:14];
  assign S1__125 = e__16[26:13] ^ e__16[31:18] ^ e__16[13:0];
  assign S1__124 = e__16[12:6] ^ e__16[17:11] ^ e__16[31:25];
  assign s_0__1 = {s_0__51, s_0__50, s_0__49, s_0__48};
  assign s_1__1 = {s_1__51, s_1__50, s_1__49, s_1__48};
  assign S0__111 = a__12[1:0] ^ a__12[12:11] ^ a__12[21:20];
  assign S0__110 = a__12[31:21] ^ a__12[10:0] ^ a__12[19:9];
  assign S0__109 = a__12[20:12] ^ a__12[31:23] ^ a__12[8:0];
  assign S0__108 = a__12[11:2] ^ a__12[22:13] ^ a__12[31:22];
  assign and_57349 = a__12 & a__11;
  assign S1__16 = {S1__127, S1__126, S1__125, S1__124};
  assign value__1 = message[511:480] + s_0__1;
  assign value__2 = w_im15__8 + s_1__1;
  assign S0__12 = {S0__111, S0__110, S0__109, S0__108};
  assign maj__12 = and_57349 ^ a__12 & a__10 ^ and_57262;
  assign temp1__65 = e__13 + S1__16;
  assign ch__16 = e__16 & e__15 ^ ~(e__16 | ~e__14);
  assign value__3 = value__1 + value__2;
  assign s_0__55 = message[422:420] ^ message[433:431];
  assign s_0__54 = message[419:416] ^ message[430:427] ^ message[447:444];
  assign s_0__53 = message[447:437] ^ message[426:416] ^ message[443:433];
  assign s_0__52 = message[436:423] ^ message[447:434] ^ message[432:419];
  assign s_1__55 = message[16:7] ^ message[18:9];
  assign s_1__54 = message[6:0] ^ message[8:2] ^ message[31:25];
  assign s_1__53 = message[31:30] ^ message[1:0] ^ message[24:23];
  assign s_1__52 = message[29:17] ^ message[31:19] ^ message[22:10];
  assign temp2__12 = S0__12 + maj__12;
  assign temp1__66 = temp1__65 + ch__16;
  assign temp1__274 = value__3 + 32'he49b_69c1;
  assign w_init_im15 = message[479:448];
  assign s_0__2 = {s_0__55, s_0__54, s_0__53, s_0__52};
  assign w_im15__9 = message[191:160];
  assign s_1__2 = {s_1__55, s_1__54, s_1__53, s_1__52};
  assign a__13 = temp1__430 + temp2__12;
  assign temp1__68 = temp1__66 + temp1__274;
  assign value__4 = w_init_im15 + s_0__2;
  assign value__5 = w_im15__9 + s_1__2;
  assign e__17 = a__13 + temp1__68;
  assign value__6 = value__4 + value__5;
  assign S0__115 = a__13[1:0] ^ a__13[12:11] ^ a__13[21:20];
  assign S0__114 = a__13[31:21] ^ a__13[10:0] ^ a__13[19:9];
  assign S0__113 = a__13[20:12] ^ a__13[31:23] ^ a__13[8:0];
  assign S0__112 = a__13[11:2] ^ a__13[22:13] ^ a__13[31:22];
  assign and_57435 = a__13 & a__12;
  assign S1__131 = e__17[5:0] ^ e__17[10:5] ^ e__17[24:19];
  assign S1__130 = e__17[31:27] ^ e__17[4:0] ^ e__17[18:14];
  assign S1__129 = e__17[26:13] ^ e__17[31:18] ^ e__17[13:0];
  assign S1__128 = e__17[12:6] ^ e__17[17:11] ^ e__17[31:25];
  assign add_57443 = value__6[31:1] + 31'h77df_23c3;
  assign S0__13 = {S0__115, S0__114, S0__113, S0__112};
  assign maj__13 = and_57435 ^ a__13 & a__11 ^ and_57349;
  assign S1__17 = {S1__131, S1__130, S1__129, S1__128};
  assign ch__17 = e__17 & e__16 ^ ~(e__17 | ~e__15);
  assign temp1__275 = {add_57443, value__6[0]};
  assign s_0__59 = message[390:388] ^ message[401:399];
  assign s_0__58 = message[387:384] ^ message[398:395] ^ message[415:412];
  assign s_0__57 = message[415:405] ^ message[394:384] ^ message[411:401];
  assign s_0__56 = message[404:391] ^ message[415:402] ^ message[400:387];
  assign s_1__59 = value__3[16:7] ^ value__3[18:9];
  assign s_1__58 = value__3[6:0] ^ value__3[8:2] ^ value__3[31:25];
  assign s_1__57 = value__3[31:30] ^ value__3[1:0] ^ value__3[24:23];
  assign s_1__56 = value__3[29:17] ^ value__3[31:19] ^ value__3[22:10];
  assign temp2__13 = S0__13 + maj__13;
  assign temp1__419 = e__14 + S1__17;
  assign temp1__420 = ch__17 + temp1__275;
  assign s_0__3 = {s_0__59, s_0__58, s_0__57, s_0__56};
  assign s_1__3 = {s_1__59, s_1__58, s_1__57, s_1__56};
  assign a__14 = temp1__427 + temp2__13;
  assign temp1__421 = temp1__419 + temp1__420;
  assign value__7 = w_im15__1 + s_0__3;
  assign value__8 = w_im15__10 + s_1__3;
  assign e__18 = a__14 + temp1__421;
  assign value__9 = value__7 + value__8;
  assign S0__119 = a__14[1:0] ^ a__14[12:11] ^ a__14[21:20];
  assign S0__118 = a__14[31:21] ^ a__14[10:0] ^ a__14[19:9];
  assign S0__117 = a__14[20:12] ^ a__14[31:23] ^ a__14[8:0];
  assign S0__116 = a__14[11:2] ^ a__14[22:13] ^ a__14[31:22];
  assign and_57522 = a__14 & a__13;
  assign S1__135 = e__18[5:0] ^ e__18[10:5] ^ e__18[24:19];
  assign S1__134 = e__18[31:27] ^ e__18[4:0] ^ e__18[18:14];
  assign S1__133 = e__18[26:13] ^ e__18[31:18] ^ e__18[13:0];
  assign S1__132 = e__18[12:6] ^ e__18[17:11] ^ e__18[31:25];
  assign add_57530 = value__9[31:1] + 31'h07e0_cee3;
  assign S0__14 = {S0__119, S0__118, S0__117, S0__116};
  assign maj__14 = and_57522 ^ a__14 & a__12 ^ and_57435;
  assign S1__18 = {S1__135, S1__134, S1__133, S1__132};
  assign ch__18 = e__18 & e__17 ^ ~(e__18 | ~e__16);
  assign temp1__276 = {add_57530, value__9[0]};
  assign s_0__63 = message[358:356] ^ message[369:367];
  assign s_0__62 = message[355:352] ^ message[366:363] ^ message[383:380];
  assign s_0__61 = message[383:373] ^ message[362:352] ^ message[379:369];
  assign s_0__60 = message[372:359] ^ message[383:370] ^ message[368:355];
  assign s_1__63 = value__6[16:7] ^ value__6[18:9];
  assign s_1__62 = value__6[6:0] ^ value__6[8:2] ^ value__6[31:25];
  assign s_1__61 = value__6[31:30] ^ value__6[1:0] ^ value__6[24:23];
  assign s_1__60 = value__6[29:17] ^ value__6[31:19] ^ value__6[22:10];
  assign temp2__14 = S0__14 + maj__14;
  assign temp1__416 = e__15 + S1__18;
  assign temp1__417 = ch__18 + temp1__276;
  assign w_im15__2 = message[415:384];
  assign s_0__4 = {s_0__63, s_0__62, s_0__61, s_0__60};
  assign w_im15__11 = message[127:96];
  assign s_1__4 = {s_1__63, s_1__62, s_1__61, s_1__60};
  assign a__15 = temp1__60 + temp2__14;
  assign temp1__418 = temp1__416 + temp1__417;
  assign value__10 = w_im15__2 + s_0__4;
  assign value__11 = w_im15__11 + s_1__4;
  assign e__19 = a__15 + temp1__418;
  assign value__12 = value__10 + value__11;
  assign S0__123 = a__15[1:0] ^ a__15[12:11] ^ a__15[21:20];
  assign S0__122 = a__15[31:21] ^ a__15[10:0] ^ a__15[19:9];
  assign S0__121 = a__15[20:12] ^ a__15[31:23] ^ a__15[8:0];
  assign S0__120 = a__15[11:2] ^ a__15[22:13] ^ a__15[31:22];
  assign and_57611 = a__15 & a__14;
  assign S1__139 = e__19[5:0] ^ e__19[10:5] ^ e__19[24:19];
  assign S1__138 = e__19[31:27] ^ e__19[4:0] ^ e__19[18:14];
  assign S1__137 = e__19[26:13] ^ e__19[31:18] ^ e__19[13:0];
  assign S1__136 = e__19[12:6] ^ e__19[17:11] ^ e__19[31:25];
  assign add_57619 = value__12[31:2] + 30'h0903_2873;
  assign S0__15 = {S0__123, S0__122, S0__121, S0__120};
  assign maj__15 = and_57611 ^ a__15 & a__13 ^ and_57522;
  assign S1__19 = {S1__139, S1__138, S1__137, S1__136};
  assign ch__19 = e__19 & e__18 ^ ~(e__19 | ~e__17);
  assign temp1__277 = {add_57619, value__12[1:0]};
  assign temp2__15 = S0__15 + maj__15;
  assign temp1__413 = e__16 + S1__19;
  assign temp1__414 = ch__19 + temp1__277;
  assign a__16 = temp1__424 + temp2__15;
  assign temp1__415 = temp1__413 + temp1__414;
  assign e__20 = a__16 + temp1__415;
  assign s_0__67 = message[326:324] ^ message[337:335];
  assign s_0__66 = message[323:320] ^ message[334:331] ^ message[351:348];
  assign s_0__65 = message[351:341] ^ message[330:320] ^ message[347:337];
  assign s_0__64 = message[340:327] ^ message[351:338] ^ message[336:323];
  assign s_1__67 = value__9[16:7] ^ value__9[18:9];
  assign s_1__66 = value__9[6:0] ^ value__9[8:2] ^ value__9[31:25];
  assign s_1__65 = value__9[31:30] ^ value__9[1:0] ^ value__9[24:23];
  assign s_1__64 = value__9[29:17] ^ value__9[31:19] ^ value__9[22:10];
  assign S1__143 = e__20[5:0] ^ e__20[10:5] ^ e__20[24:19];
  assign S1__142 = e__20[31:27] ^ e__20[4:0] ^ e__20[18:14];
  assign S1__141 = e__20[26:13] ^ e__20[31:18] ^ e__20[13:0];
  assign S1__140 = e__20[12:6] ^ e__20[17:11] ^ e__20[31:25];
  assign s_0__5 = {s_0__67, s_0__66, s_0__65, s_0__64};
  assign w_im15__12 = message[95:64];
  assign s_1__5 = {s_1__67, s_1__66, s_1__65, s_1__64};
  assign S0__127 = a__16[1:0] ^ a__16[12:11] ^ a__16[21:20];
  assign S0__126 = a__16[31:21] ^ a__16[10:0] ^ a__16[19:9];
  assign S0__125 = a__16[20:12] ^ a__16[31:23] ^ a__16[8:0];
  assign S0__124 = a__16[11:2] ^ a__16[22:13] ^ a__16[31:22];
  assign and_57698 = a__16 & a__15;
  assign S1__20 = {S1__143, S1__142, S1__141, S1__140};
  assign value__13 = w_im15__3 + s_0__5;
  assign value__14 = w_im15__12 + s_1__5;
  assign S0__16 = {S0__127, S0__126, S0__125, S0__124};
  assign maj__16 = and_57698 ^ a__16 & a__14 ^ and_57611;
  assign temp1__81 = e__17 + S1__20;
  assign ch__20 = e__20 & e__19 ^ ~(e__20 | ~e__18);
  assign value__15 = value__13 + value__14;
  assign s_0__71 = message[294:292] ^ message[305:303];
  assign s_0__70 = message[291:288] ^ message[302:299] ^ message[319:316];
  assign s_0__69 = message[319:309] ^ message[298:288] ^ message[315:305];
  assign s_0__68 = message[308:295] ^ message[319:306] ^ message[304:291];
  assign s_1__71 = value__12[16:7] ^ value__12[18:9];
  assign s_1__70 = value__12[6:0] ^ value__12[8:2] ^ value__12[31:25];
  assign s_1__69 = value__12[31:30] ^ value__12[1:0] ^ value__12[24:23];
  assign s_1__68 = value__12[29:17] ^ value__12[31:19] ^ value__12[22:10];
  assign temp2__16 = S0__16 + maj__16;
  assign temp1__82 = temp1__81 + ch__20;
  assign temp1__278 = value__15 + 32'h2de9_2c6f;
  assign s_0__6 = {s_0__71, s_0__70, s_0__69, s_0__68};
  assign s_1__6 = {s_1__71, s_1__70, s_1__69, s_1__68};
  assign a__17 = temp1__68 + temp2__16;
  assign temp1__84 = temp1__82 + temp1__278;
  assign value__16 = w_im15__4 + s_0__6;
  assign value__17 = w_init_im2 + s_1__6;
  assign e__21 = a__17 + temp1__84;
  assign value__18 = value__16 + value__17;
  assign S0__131 = a__17[1:0] ^ a__17[12:11] ^ a__17[21:20];
  assign S0__130 = a__17[31:21] ^ a__17[10:0] ^ a__17[19:9];
  assign S0__129 = a__17[20:12] ^ a__17[31:23] ^ a__17[8:0];
  assign S0__128 = a__17[11:2] ^ a__17[22:13] ^ a__17[31:22];
  assign and_57782 = a__17 & a__16;
  assign S1__147 = e__21[5:0] ^ e__21[10:5] ^ e__21[24:19];
  assign S1__146 = e__21[31:27] ^ e__21[4:0] ^ e__21[18:14];
  assign S1__145 = e__21[26:13] ^ e__21[31:18] ^ e__21[13:0];
  assign S1__144 = e__21[12:6] ^ e__21[17:11] ^ e__21[31:25];
  assign add_57790 = value__18[31:1] + 31'h253a_4255;
  assign S0__17 = {S0__131, S0__130, S0__129, S0__128};
  assign maj__17 = and_57782 ^ a__17 & a__15 ^ and_57698;
  assign S1__21 = {S1__147, S1__146, S1__145, S1__144};
  assign ch__21 = e__21 & e__20 ^ ~(e__21 | ~e__19);
  assign temp1__279 = {add_57790, value__18[0]};
  assign s_0__75 = message[262:260] ^ message[273:271];
  assign s_0__74 = message[259:256] ^ message[270:267] ^ message[287:284];
  assign s_0__73 = message[287:277] ^ message[266:256] ^ message[283:273];
  assign s_0__72 = message[276:263] ^ message[287:274] ^ message[272:259];
  assign s_1__75 = value__15[16:7] ^ value__15[18:9];
  assign s_1__74 = value__15[6:0] ^ value__15[8:2] ^ value__15[31:25];
  assign s_1__73 = value__15[31:30] ^ value__15[1:0] ^ value__15[24:23];
  assign s_1__72 = value__15[29:17] ^ value__15[31:19] ^ value__15[22:10];
  assign temp2__17 = S0__17 + maj__17;
  assign temp1__410 = e__18 + S1__21;
  assign temp1__411 = ch__21 + temp1__279;
  assign w_im15__5 = message[319:288];
  assign s_0__7 = {s_0__75, s_0__74, s_0__73, s_0__72};
  assign w_im2__1 = message[31:0];
  assign s_1__7 = {s_1__75, s_1__74, s_1__73, s_1__72};
  assign a__18 = temp1__421 + temp2__17;
  assign temp1__412 = temp1__410 + temp1__411;
  assign value__19 = w_im15__5 + s_0__7;
  assign value__20 = w_im2__1 + s_1__7;
  assign e__22 = a__18 + temp1__412;
  assign value__21 = value__19 + value__20;
  assign S0__135 = a__18[1:0] ^ a__18[12:11] ^ a__18[21:20];
  assign S0__134 = a__18[31:21] ^ a__18[10:0] ^ a__18[19:9];
  assign S0__133 = a__18[20:12] ^ a__18[31:23] ^ a__18[8:0];
  assign S0__132 = a__18[11:2] ^ a__18[22:13] ^ a__18[31:22];
  assign and_57871 = a__18 & a__17;
  assign S1__151 = e__22[5:0] ^ e__22[10:5] ^ e__22[24:19];
  assign S1__150 = e__22[31:27] ^ e__22[4:0] ^ e__22[18:14];
  assign S1__149 = e__22[26:13] ^ e__22[31:18] ^ e__22[13:0];
  assign S1__148 = e__22[12:6] ^ e__22[17:11] ^ e__22[31:25];
  assign add_57879 = value__21[31:2] + 30'h172c_2a77;
  assign S0__18 = {S0__135, S0__134, S0__133, S0__132};
  assign maj__18 = and_57871 ^ a__18 & a__16 ^ and_57782;
  assign S1__22 = {S1__151, S1__150, S1__149, S1__148};
  assign ch__22 = e__22 & e__21 ^ ~(e__22 | ~e__20);
  assign temp1__280 = {add_57879, value__21[1:0]};
  assign s_0__79 = message[230:228] ^ message[241:239];
  assign s_0__78 = message[227:224] ^ message[238:235] ^ message[255:252];
  assign s_0__77 = message[255:245] ^ message[234:224] ^ message[251:241];
  assign s_0__76 = message[244:231] ^ message[255:242] ^ message[240:227];
  assign s_1__79 = value__18[16:7] ^ value__18[18:9];
  assign s_1__78 = value__18[6:0] ^ value__18[8:2] ^ value__18[31:25];
  assign s_1__77 = value__18[31:30] ^ value__18[1:0] ^ value__18[24:23];
  assign s_1__76 = value__18[29:17] ^ value__18[31:19] ^ value__18[22:10];
  assign temp2__18 = S0__18 + maj__18;
  assign temp1__407 = e__19 + S1__22;
  assign temp1__408 = ch__22 + temp1__280;
  assign s_0__8 = {s_0__79, s_0__78, s_0__77, s_0__76};
  assign s_1__8 = {s_1__79, s_1__78, s_1__77, s_1__76};
  assign a__19 = temp1__418 + temp2__18;
  assign temp1__409 = temp1__407 + temp1__408;
  assign value__22 = w_im15__6 + s_0__8;
  assign value__23 = value__3 + s_1__8;
  assign e__23 = a__19 + temp1__409;
  assign value__24 = value__22 + value__23;
  assign S0__139 = a__19[1:0] ^ a__19[12:11] ^ a__19[21:20];
  assign S0__138 = a__19[31:21] ^ a__19[10:0] ^ a__19[19:9];
  assign S0__137 = a__19[20:12] ^ a__19[31:23] ^ a__19[8:0];
  assign S0__136 = a__19[11:2] ^ a__19[22:13] ^ a__19[31:22];
  assign and_57958 = a__19 & a__18;
  assign S1__155 = e__23[5:0] ^ e__23[10:5] ^ e__23[24:19];
  assign S1__154 = e__23[31:27] ^ e__23[4:0] ^ e__23[18:14];
  assign S1__153 = e__23[26:13] ^ e__23[31:18] ^ e__23[13:0];
  assign S1__152 = e__23[12:6] ^ e__23[17:11] ^ e__23[31:25];
  assign add_57966 = value__24[31:1] + 31'h3b7c_c46d;
  assign S0__19 = {S0__139, S0__138, S0__137, S0__136};
  assign maj__19 = and_57958 ^ a__19 & a__17 ^ and_57871;
  assign S1__23 = {S1__155, S1__154, S1__153, S1__152};
  assign ch__23 = e__23 & e__22 ^ ~(e__23 | ~e__21);
  assign temp1__281 = {add_57966, value__24[0]};
  assign s_0__83 = message[198:196] ^ message[209:207];
  assign s_0__82 = message[195:192] ^ message[206:203] ^ message[223:220];
  assign s_0__81 = message[223:213] ^ message[202:192] ^ message[219:209];
  assign s_0__80 = message[212:199] ^ message[223:210] ^ message[208:195];
  assign s_1__83 = value__21[16:7] ^ value__21[18:9];
  assign s_1__82 = value__21[6:0] ^ value__21[8:2] ^ value__21[31:25];
  assign s_1__81 = value__21[31:30] ^ value__21[1:0] ^ value__21[24:23];
  assign s_1__80 = value__21[29:17] ^ value__21[31:19] ^ value__21[22:10];
  assign temp2__19 = S0__19 + maj__19;
  assign temp1__404 = e__20 + S1__23;
  assign temp1__405 = ch__23 + temp1__281;
  assign w_im15__7 = message[255:224];
  assign s_0__9 = {s_0__83, s_0__82, s_0__81, s_0__80};
  assign s_1__9 = {s_1__83, s_1__82, s_1__81, s_1__80};
  assign a__20 = temp1__415 + temp2__19;
  assign temp1__406 = temp1__404 + temp1__405;
  assign value__25 = w_im15__7 + s_0__9;
  assign value__26 = value__6 + s_1__9;
  assign e__24 = a__20 + temp1__406;
  assign value__27 = value__25 + value__26;
  assign S0__143 = a__20[1:0] ^ a__20[12:11] ^ a__20[21:20];
  assign S0__142 = a__20[31:21] ^ a__20[10:0] ^ a__20[19:9];
  assign S0__141 = a__20[20:12] ^ a__20[31:23] ^ a__20[8:0];
  assign S0__140 = a__20[11:2] ^ a__20[22:13] ^ a__20[31:22];
  assign and_58045 = a__20 & a__19;
  assign S1__159 = e__24[5:0] ^ e__24[10:5] ^ e__24[24:19];
  assign S1__158 = e__24[31:27] ^ e__24[4:0] ^ e__24[18:14];
  assign S1__157 = e__24[26:13] ^ e__24[31:18] ^ e__24[13:0];
  assign S1__156 = e__24[12:6] ^ e__24[17:11] ^ e__24[31:25];
  assign add_58053 = value__27[31:1] + 31'h4c1f_28a9;
  assign S0__20 = {S0__143, S0__142, S0__141, S0__140};
  assign maj__20 = and_58045 ^ a__20 & a__18 ^ and_57958;
  assign S1__24 = {S1__159, S1__158, S1__157, S1__156};
  assign ch__24 = e__24 & e__23 ^ ~(e__24 | ~e__22);
  assign temp1__282 = {add_58053, value__27[0]};
  assign temp2__20 = S0__20 + maj__20;
  assign temp1__401 = e__21 + S1__24;
  assign temp1__402 = ch__24 + temp1__282;
  assign a__21 = temp1__84 + temp2__20;
  assign temp1__403 = temp1__401 + temp1__402;
  assign e__25 = a__21 + temp1__403;
  assign s_0__87 = message[166:164] ^ message[177:175];
  assign s_0__86 = message[163:160] ^ message[174:171] ^ message[191:188];
  assign s_0__85 = message[191:181] ^ message[170:160] ^ message[187:177];
  assign s_0__84 = message[180:167] ^ message[191:178] ^ message[176:163];
  assign s_1__87 = value__24[16:7] ^ value__24[18:9];
  assign s_1__86 = value__24[6:0] ^ value__24[8:2] ^ value__24[31:25];
  assign s_1__85 = value__24[31:30] ^ value__24[1:0] ^ value__24[24:23];
  assign s_1__84 = value__24[29:17] ^ value__24[31:19] ^ value__24[22:10];
  assign S1__163 = e__25[5:0] ^ e__25[10:5] ^ e__25[24:19];
  assign S1__162 = e__25[31:27] ^ e__25[4:0] ^ e__25[18:14];
  assign S1__161 = e__25[26:13] ^ e__25[31:18] ^ e__25[13:0];
  assign S1__160 = e__25[12:6] ^ e__25[17:11] ^ e__25[31:25];
  assign s_0__10 = {s_0__87, s_0__86, s_0__85, s_0__84};
  assign s_1__10 = {s_1__87, s_1__86, s_1__85, s_1__84};
  assign S0__147 = a__21[1:0] ^ a__21[12:11] ^ a__21[21:20];
  assign S0__146 = a__21[31:21] ^ a__21[10:0] ^ a__21[19:9];
  assign S0__145 = a__21[20:12] ^ a__21[31:23] ^ a__21[8:0];
  assign S0__144 = a__21[11:2] ^ a__21[22:13] ^ a__21[31:22];
  assign and_58131 = a__21 & a__20;
  assign S1__25 = {S1__163, S1__162, S1__161, S1__160};
  assign value__28 = w_im15__8 + s_0__10;
  assign value__29 = value__9 + s_1__10;
  assign S0__21 = {S0__147, S0__146, S0__145, S0__144};
  assign maj__21 = and_58131 ^ a__21 & a__19 ^ and_58045;
  assign temp1__101 = e__22 + S1__25;
  assign ch__25 = e__25 & e__24 ^ ~(e__25 | ~e__23);
  assign value__30 = value__28 + value__29;
  assign s_0__91 = message[134:132] ^ message[145:143];
  assign s_0__90 = message[131:128] ^ message[142:139] ^ message[159:156];
  assign s_0__89 = message[159:149] ^ message[138:128] ^ message[155:145];
  assign s_0__88 = message[148:135] ^ message[159:146] ^ message[144:131];
  assign s_1__91 = value__27[16:7] ^ value__27[18:9];
  assign s_1__90 = value__27[6:0] ^ value__27[8:2] ^ value__27[31:25];
  assign s_1__89 = value__27[31:30] ^ value__27[1:0] ^ value__27[24:23];
  assign s_1__88 = value__27[29:17] ^ value__27[31:19] ^ value__27[22:10];
  assign temp2__21 = S0__21 + maj__21;
  assign temp1__102 = temp1__101 + ch__25;
  assign temp1__283 = value__30 + 32'ha831_c66d;
  assign s_0__11 = {s_0__91, s_0__90, s_0__89, s_0__88};
  assign s_1__11 = {s_1__91, s_1__90, s_1__89, s_1__88};
  assign a__22 = temp1__412 + temp2__21;
  assign temp1__104 = temp1__102 + temp1__283;
  assign value__31 = w_im15__9 + s_0__11;
  assign value__32 = value__12 + s_1__11;
  assign e__26 = a__22 + temp1__104;
  assign value__33 = value__31 + value__32;
  assign S0__151 = a__22[1:0] ^ a__22[12:11] ^ a__22[21:20];
  assign S0__150 = a__22[31:21] ^ a__22[10:0] ^ a__22[19:9];
  assign S0__149 = a__22[20:12] ^ a__22[31:23] ^ a__22[8:0];
  assign S0__148 = a__22[11:2] ^ a__22[22:13] ^ a__22[31:22];
  assign and_58216 = a__22 & a__21;
  assign S1__167 = e__26[5:0] ^ e__26[10:5] ^ e__26[24:19];
  assign S1__166 = e__26[31:27] ^ e__26[4:0] ^ e__26[18:14];
  assign S1__165 = e__26[26:13] ^ e__26[31:18] ^ e__26[13:0];
  assign S1__164 = e__26[12:6] ^ e__26[17:11] ^ e__26[31:25];
  assign add_58224 = value__33[31:3] + 29'h1600_64f9;
  assign S0__22 = {S0__151, S0__150, S0__149, S0__148};
  assign maj__22 = and_58216 ^ a__22 & a__20 ^ and_58131;
  assign S1__26 = {S1__167, S1__166, S1__165, S1__164};
  assign ch__26 = e__26 & e__25 ^ ~(e__26 | ~e__24);
  assign temp1__284 = {add_58224, value__33[2:0]};
  assign temp2__22 = S0__22 + maj__22;
  assign temp1__398 = e__23 + S1__26;
  assign temp1__399 = ch__26 + temp1__284;
  assign a__23 = temp1__409 + temp2__22;
  assign temp1__400 = temp1__398 + temp1__399;
  assign e__27 = a__23 + temp1__400;
  assign s_0__95 = message[102:100] ^ message[113:111];
  assign s_0__94 = message[99:96] ^ message[110:107] ^ message[127:124];
  assign s_0__93 = message[127:117] ^ message[106:96] ^ message[123:113];
  assign s_0__92 = message[116:103] ^ message[127:114] ^ message[112:99];
  assign s_1__95 = value__30[16:7] ^ value__30[18:9];
  assign s_1__94 = value__30[6:0] ^ value__30[8:2] ^ value__30[31:25];
  assign s_1__93 = value__30[31:30] ^ value__30[1:0] ^ value__30[24:23];
  assign s_1__92 = value__30[29:17] ^ value__30[31:19] ^ value__30[22:10];
  assign S1__171 = e__27[5:0] ^ e__27[10:5] ^ e__27[24:19];
  assign S1__170 = e__27[31:27] ^ e__27[4:0] ^ e__27[18:14];
  assign S1__169 = e__27[26:13] ^ e__27[31:18] ^ e__27[13:0];
  assign S1__168 = e__27[12:6] ^ e__27[17:11] ^ e__27[31:25];
  assign s_0__12 = {s_0__95, s_0__94, s_0__93, s_0__92};
  assign s_1__12 = {s_1__95, s_1__94, s_1__93, s_1__92};
  assign S0__155 = a__23[1:0] ^ a__23[12:11] ^ a__23[21:20];
  assign S0__154 = a__23[31:21] ^ a__23[10:0] ^ a__23[19:9];
  assign S0__153 = a__23[20:12] ^ a__23[31:23] ^ a__23[8:0];
  assign S0__152 = a__23[11:2] ^ a__23[22:13] ^ a__23[31:22];
  assign and_58302 = a__23 & a__22;
  assign S1__27 = {S1__171, S1__170, S1__169, S1__168};
  assign value__34 = w_im15__10 + s_0__12;
  assign value__35 = value__15 + s_1__12;
  assign S0__23 = {S0__155, S0__154, S0__153, S0__152};
  assign maj__23 = and_58302 ^ a__23 & a__21 ^ and_58216;
  assign temp1__109 = e__24 + S1__27;
  assign ch__27 = e__27 & e__26 ^ ~(e__27 | ~e__25);
  assign value__36 = value__34 + value__35;
  assign temp2__23 = S0__23 + maj__23;
  assign temp1__110 = temp1__109 + ch__27;
  assign temp1__285 = value__36 + 32'hbf59_7fc7;
  assign a__24 = temp1__406 + temp2__23;
  assign temp1__112 = temp1__110 + temp1__285;
  assign e__28 = a__24 + temp1__112;
  assign s_0__99 = message[70:68] ^ message[81:79];
  assign s_0__98 = message[67:64] ^ message[78:75] ^ message[95:92];
  assign s_0__97 = message[95:85] ^ message[74:64] ^ message[91:81];
  assign s_0__96 = message[84:71] ^ message[95:82] ^ message[80:67];
  assign s_1__99 = value__33[16:7] ^ value__33[18:9];
  assign s_1__98 = value__33[6:0] ^ value__33[8:2] ^ value__33[31:25];
  assign s_1__97 = value__33[31:30] ^ value__33[1:0] ^ value__33[24:23];
  assign s_1__96 = value__33[29:17] ^ value__33[31:19] ^ value__33[22:10];
  assign S1__175 = e__28[5:0] ^ e__28[10:5] ^ e__28[24:19];
  assign S1__174 = e__28[31:27] ^ e__28[4:0] ^ e__28[18:14];
  assign S1__173 = e__28[26:13] ^ e__28[31:18] ^ e__28[13:0];
  assign S1__172 = e__28[12:6] ^ e__28[17:11] ^ e__28[31:25];
  assign s_0__13 = {s_0__99, s_0__98, s_0__97, s_0__96};
  assign s_1__13 = {s_1__99, s_1__98, s_1__97, s_1__96};
  assign S0__159 = a__24[1:0] ^ a__24[12:11] ^ a__24[21:20];
  assign S0__158 = a__24[31:21] ^ a__24[10:0] ^ a__24[19:9];
  assign S0__157 = a__24[20:12] ^ a__24[31:23] ^ a__24[8:0];
  assign S0__156 = a__24[11:2] ^ a__24[22:13] ^ a__24[31:22];
  assign and_58386 = a__24 & a__23;
  assign S1__28 = {S1__175, S1__174, S1__173, S1__172};
  assign value__37 = w_im15__11 + s_0__13;
  assign value__38 = value__18 + s_1__13;
  assign S0__24 = {S0__159, S0__158, S0__157, S0__156};
  assign maj__24 = and_58386 ^ a__24 & a__22 ^ and_58302;
  assign temp1__113 = e__25 + S1__28;
  assign ch__28 = e__28 & e__27 ^ ~(e__28 | ~e__26);
  assign value__39 = value__37 + value__38;
  assign temp2__24 = S0__24 + maj__24;
  assign temp1__114 = temp1__113 + ch__28;
  assign temp1__286 = value__39 + 32'hc6e0_0bf3;
  assign a__25 = temp1__403 + temp2__24;
  assign temp1__116 = temp1__114 + temp1__286;
  assign e__29 = a__25 + temp1__116;
  assign s_0__103 = message[38:36] ^ message[49:47];
  assign s_0__102 = message[35:32] ^ message[46:43] ^ message[63:60];
  assign s_0__101 = message[63:53] ^ message[42:32] ^ message[59:49];
  assign s_0__100 = message[52:39] ^ message[63:50] ^ message[48:35];
  assign s_1__103 = value__36[16:7] ^ value__36[18:9];
  assign s_1__102 = value__36[6:0] ^ value__36[8:2] ^ value__36[31:25];
  assign s_1__101 = value__36[31:30] ^ value__36[1:0] ^ value__36[24:23];
  assign s_1__100 = value__36[29:17] ^ value__36[31:19] ^ value__36[22:10];
  assign S1__179 = e__29[5:0] ^ e__29[10:5] ^ e__29[24:19];
  assign S1__178 = e__29[31:27] ^ e__29[4:0] ^ e__29[18:14];
  assign S1__177 = e__29[26:13] ^ e__29[31:18] ^ e__29[13:0];
  assign S1__176 = e__29[12:6] ^ e__29[17:11] ^ e__29[31:25];
  assign s_0__14 = {s_0__103, s_0__102, s_0__101, s_0__100};
  assign s_1__14 = {s_1__103, s_1__102, s_1__101, s_1__100};
  assign S0__163 = a__25[1:0] ^ a__25[12:11] ^ a__25[21:20];
  assign S0__162 = a__25[31:21] ^ a__25[10:0] ^ a__25[19:9];
  assign S0__161 = a__25[20:12] ^ a__25[31:23] ^ a__25[8:0];
  assign S0__160 = a__25[11:2] ^ a__25[22:13] ^ a__25[31:22];
  assign and_58470 = a__25 & a__24;
  assign S1__29 = {S1__179, S1__178, S1__177, S1__176};
  assign value__40 = w_im15__12 + s_0__14;
  assign value__41 = value__21 + s_1__14;
  assign S0__25 = {S0__163, S0__162, S0__161, S0__160};
  assign maj__25 = and_58470 ^ a__25 & a__23 ^ and_58386;
  assign temp1__117 = e__26 + S1__29;
  assign ch__29 = e__29 & e__28 ^ ~(e__29 | ~e__27);
  assign value__42 = value__40 + value__41;
  assign temp2__25 = S0__25 + maj__25;
  assign temp1__118 = temp1__117 + ch__29;
  assign temp1__287 = value__42 + 32'hd5a7_9147;
  assign a__26 = temp1__104 + temp2__25;
  assign temp1__120 = temp1__118 + temp1__287;
  assign e__30 = a__26 + temp1__120;
  assign s_0__107 = message[6:4] ^ message[17:15];
  assign s_0__106 = message[3:0] ^ message[14:11] ^ message[31:28];
  assign s_0__105 = message[31:21] ^ message[10:0] ^ message[27:17];
  assign s_0__104 = message[20:7] ^ message[31:18] ^ message[16:3];
  assign s_1__107 = value__39[16:7] ^ value__39[18:9];
  assign s_1__106 = value__39[6:0] ^ value__39[8:2] ^ value__39[31:25];
  assign s_1__105 = value__39[31:30] ^ value__39[1:0] ^ value__39[24:23];
  assign s_1__104 = value__39[29:17] ^ value__39[31:19] ^ value__39[22:10];
  assign S1__183 = e__30[5:0] ^ e__30[10:5] ^ e__30[24:19];
  assign S1__182 = e__30[31:27] ^ e__30[4:0] ^ e__30[18:14];
  assign S1__181 = e__30[26:13] ^ e__30[31:18] ^ e__30[13:0];
  assign S1__180 = e__30[12:6] ^ e__30[17:11] ^ e__30[31:25];
  assign s_0__15 = {s_0__107, s_0__106, s_0__105, s_0__104};
  assign s_1__15 = {s_1__107, s_1__106, s_1__105, s_1__104};
  assign S0__167 = a__26[1:0] ^ a__26[12:11] ^ a__26[21:20];
  assign S0__166 = a__26[31:21] ^ a__26[10:0] ^ a__26[19:9];
  assign S0__165 = a__26[20:12] ^ a__26[31:23] ^ a__26[8:0];
  assign S0__164 = a__26[11:2] ^ a__26[22:13] ^ a__26[31:22];
  assign and_58554 = a__26 & a__25;
  assign S1__30 = {S1__183, S1__182, S1__181, S1__180};
  assign value__43 = w_init_im2 + s_0__15;
  assign value__44 = value__24 + s_1__15;
  assign S0__26 = {S0__167, S0__166, S0__165, S0__164};
  assign maj__26 = and_58554 ^ a__26 & a__24 ^ and_58470;
  assign temp1__121 = e__27 + S1__30;
  assign ch__30 = e__30 & e__29 ^ ~(e__30 | ~e__28);
  assign value__45 = value__43 + value__44;
  assign temp2__26 = S0__26 + maj__26;
  assign temp1__122 = temp1__121 + ch__30;
  assign temp1__288 = value__45 + 32'h06ca_6351;
  assign a__27 = temp1__400 + temp2__26;
  assign temp1__124 = temp1__122 + temp1__288;
  assign e__31 = a__27 + temp1__124;
  assign s_0__111 = value__3[6:4] ^ value__3[17:15];
  assign s_0__110 = value__3[3:0] ^ value__3[14:11] ^ value__3[31:28];
  assign s_0__109 = value__3[31:21] ^ value__3[10:0] ^ value__3[27:17];
  assign s_0__108 = value__3[20:7] ^ value__3[31:18] ^ value__3[16:3];
  assign s_1__111 = value__42[16:7] ^ value__42[18:9];
  assign s_1__110 = value__42[6:0] ^ value__42[8:2] ^ value__42[31:25];
  assign s_1__109 = value__42[31:30] ^ value__42[1:0] ^ value__42[24:23];
  assign s_1__108 = value__42[29:17] ^ value__42[31:19] ^ value__42[22:10];
  assign S1__187 = e__31[5:0] ^ e__31[10:5] ^ e__31[24:19];
  assign S1__186 = e__31[31:27] ^ e__31[4:0] ^ e__31[18:14];
  assign S1__185 = e__31[26:13] ^ e__31[31:18] ^ e__31[13:0];
  assign S1__184 = e__31[12:6] ^ e__31[17:11] ^ e__31[31:25];
  assign s_0__16 = {s_0__111, s_0__110, s_0__109, s_0__108};
  assign s_1__16 = {s_1__111, s_1__110, s_1__109, s_1__108};
  assign S0__171 = a__27[1:0] ^ a__27[12:11] ^ a__27[21:20];
  assign S0__170 = a__27[31:21] ^ a__27[10:0] ^ a__27[19:9];
  assign S0__169 = a__27[20:12] ^ a__27[31:23] ^ a__27[8:0];
  assign S0__168 = a__27[11:2] ^ a__27[22:13] ^ a__27[31:22];
  assign and_58638 = a__27 & a__26;
  assign S1__31 = {S1__187, S1__186, S1__185, S1__184};
  assign value__46 = w_im2__1 + s_0__16;
  assign value__47 = value__27 + s_1__16;
  assign S0__27 = {S0__171, S0__170, S0__169, S0__168};
  assign maj__27 = and_58638 ^ a__27 & a__25 ^ and_58554;
  assign temp1__125 = e__28 + S1__31;
  assign ch__31 = e__31 & e__30 ^ ~(e__31 | ~e__29);
  assign value__48 = value__46 + value__47;
  assign temp2__27 = S0__27 + maj__27;
  assign temp1__126 = temp1__125 + ch__31;
  assign temp1__289 = value__48 + 32'h1429_2967;
  assign a__28 = temp1__112 + temp2__27;
  assign temp1__128 = temp1__126 + temp1__289;
  assign e__32 = a__28 + temp1__128;
  assign s_0__115 = value__6[6:4] ^ value__6[17:15];
  assign s_0__114 = value__6[3:0] ^ value__6[14:11] ^ value__6[31:28];
  assign s_0__113 = value__6[31:21] ^ value__6[10:0] ^ value__6[27:17];
  assign s_0__112 = value__6[20:7] ^ value__6[31:18] ^ value__6[16:3];
  assign s_1__115 = value__45[16:7] ^ value__45[18:9];
  assign s_1__114 = value__45[6:0] ^ value__45[8:2] ^ value__45[31:25];
  assign s_1__113 = value__45[31:30] ^ value__45[1:0] ^ value__45[24:23];
  assign s_1__112 = value__45[29:17] ^ value__45[31:19] ^ value__45[22:10];
  assign S1__191 = e__32[5:0] ^ e__32[10:5] ^ e__32[24:19];
  assign S1__190 = e__32[31:27] ^ e__32[4:0] ^ e__32[18:14];
  assign S1__189 = e__32[26:13] ^ e__32[31:18] ^ e__32[13:0];
  assign S1__188 = e__32[12:6] ^ e__32[17:11] ^ e__32[31:25];
  assign s_0__17 = {s_0__115, s_0__114, s_0__113, s_0__112};
  assign s_1__17 = {s_1__115, s_1__114, s_1__113, s_1__112};
  assign S0__175 = a__28[1:0] ^ a__28[12:11] ^ a__28[21:20];
  assign S0__174 = a__28[31:21] ^ a__28[10:0] ^ a__28[19:9];
  assign S0__173 = a__28[20:12] ^ a__28[31:23] ^ a__28[8:0];
  assign S0__172 = a__28[11:2] ^ a__28[22:13] ^ a__28[31:22];
  assign and_58722 = a__28 & a__27;
  assign S1__32 = {S1__191, S1__190, S1__189, S1__188};
  assign value__49 = value__3 + s_0__17;
  assign value__50 = value__30 + s_1__17;
  assign S0__28 = {S0__175, S0__174, S0__173, S0__172};
  assign maj__28 = and_58722 ^ a__28 & a__26 ^ and_58638;
  assign temp1__129 = e__29 + S1__32;
  assign ch__32 = e__32 & e__31 ^ ~(e__32 | ~e__30);
  assign value__51 = value__49 + value__50;
  assign s_0__119 = value__9[6:4] ^ value__9[17:15];
  assign s_0__118 = value__9[3:0] ^ value__9[14:11] ^ value__9[31:28];
  assign s_0__117 = value__9[31:21] ^ value__9[10:0] ^ value__9[27:17];
  assign s_0__116 = value__9[20:7] ^ value__9[31:18] ^ value__9[16:3];
  assign s_1__119 = value__48[16:7] ^ value__48[18:9];
  assign s_1__118 = value__48[6:0] ^ value__48[8:2] ^ value__48[31:25];
  assign s_1__117 = value__48[31:30] ^ value__48[1:0] ^ value__48[24:23];
  assign s_1__116 = value__48[29:17] ^ value__48[31:19] ^ value__48[22:10];
  assign temp2__28 = S0__28 + maj__28;
  assign temp1__130 = temp1__129 + ch__32;
  assign temp1__290 = value__51 + 32'h27b7_0a85;
  assign s_0__18 = {s_0__119, s_0__118, s_0__117, s_0__116};
  assign s_1__18 = {s_1__119, s_1__118, s_1__117, s_1__116};
  assign a__29 = temp1__116 + temp2__28;
  assign temp1__132 = temp1__130 + temp1__290;
  assign value__52 = value__6 + s_0__18;
  assign value__53 = value__33 + s_1__18;
  assign e__33 = a__29 + temp1__132;
  assign value__54 = value__52 + value__53;
  assign S0__179 = a__29[1:0] ^ a__29[12:11] ^ a__29[21:20];
  assign S0__178 = a__29[31:21] ^ a__29[10:0] ^ a__29[19:9];
  assign S0__177 = a__29[20:12] ^ a__29[31:23] ^ a__29[8:0];
  assign S0__176 = a__29[11:2] ^ a__29[22:13] ^ a__29[31:22];
  assign and_58807 = a__29 & a__28;
  assign S1__195 = e__33[5:0] ^ e__33[10:5] ^ e__33[24:19];
  assign S1__194 = e__33[31:27] ^ e__33[4:0] ^ e__33[18:14];
  assign S1__193 = e__33[26:13] ^ e__33[31:18] ^ e__33[13:0];
  assign S1__192 = e__33[12:6] ^ e__33[17:11] ^ e__33[31:25];
  assign add_58815 = value__54[31:3] + 29'h05c3_6427;
  assign S0__29 = {S0__179, S0__178, S0__177, S0__176};
  assign maj__29 = and_58807 ^ a__29 & a__27 ^ and_58722;
  assign S1__33 = {S1__195, S1__194, S1__193, S1__192};
  assign ch__33 = e__33 & e__32 ^ ~(e__33 | ~e__31);
  assign temp1__291 = {add_58815, value__54[2:0]};
  assign s_0__123 = value__12[6:4] ^ value__12[17:15];
  assign s_0__122 = value__12[3:0] ^ value__12[14:11] ^ value__12[31:28];
  assign s_0__121 = value__12[31:21] ^ value__12[10:0] ^ value__12[27:17];
  assign s_0__120 = value__12[20:7] ^ value__12[31:18] ^ value__12[16:3];
  assign s_1__123 = value__51[16:7] ^ value__51[18:9];
  assign s_1__122 = value__51[6:0] ^ value__51[8:2] ^ value__51[31:25];
  assign s_1__121 = value__51[31:30] ^ value__51[1:0] ^ value__51[24:23];
  assign s_1__120 = value__51[29:17] ^ value__51[31:19] ^ value__51[22:10];
  assign temp2__29 = S0__29 + maj__29;
  assign temp1__395 = e__30 + S1__33;
  assign temp1__396 = ch__33 + temp1__291;
  assign s_0__19 = {s_0__123, s_0__122, s_0__121, s_0__120};
  assign s_1__19 = {s_1__123, s_1__122, s_1__121, s_1__120};
  assign a__30 = temp1__120 + temp2__29;
  assign temp1__397 = temp1__395 + temp1__396;
  assign value__55 = value__9 + s_0__19;
  assign value__56 = value__36 + s_1__19;
  assign e__34 = a__30 + temp1__397;
  assign value__57 = value__55 + value__56;
  assign S0__183 = a__30[1:0] ^ a__30[12:11] ^ a__30[21:20];
  assign S0__182 = a__30[31:21] ^ a__30[10:0] ^ a__30[19:9];
  assign S0__181 = a__30[20:12] ^ a__30[31:23] ^ a__30[8:0];
  assign S0__180 = a__30[11:2] ^ a__30[22:13] ^ a__30[31:22];
  assign and_58894 = a__30 & a__29;
  assign S1__199 = e__34[5:0] ^ e__34[10:5] ^ e__34[24:19];
  assign S1__198 = e__34[31:27] ^ e__34[4:0] ^ e__34[18:14];
  assign S1__197 = e__34[26:13] ^ e__34[31:18] ^ e__34[13:0];
  assign S1__196 = e__34[12:6] ^ e__34[17:11] ^ e__34[31:25];
  assign add_58902 = value__57[31:2] + 30'h134b_1b7f;
  assign S0__30 = {S0__183, S0__182, S0__181, S0__180};
  assign maj__30 = and_58894 ^ a__30 & a__28 ^ and_58807;
  assign S1__34 = {S1__199, S1__198, S1__197, S1__196};
  assign ch__34 = e__34 & e__33 ^ ~(e__34 | ~e__32);
  assign temp1__292 = {add_58902, value__57[1:0]};
  assign temp2__30 = S0__30 + maj__30;
  assign temp1__392 = e__31 + S1__34;
  assign temp1__393 = ch__34 + temp1__292;
  assign a__31 = temp1__124 + temp2__30;
  assign temp1__394 = temp1__392 + temp1__393;
  assign e__35 = a__31 + temp1__394;
  assign s_0__127 = value__15[6:4] ^ value__15[17:15];
  assign s_0__126 = value__15[3:0] ^ value__15[14:11] ^ value__15[31:28];
  assign s_0__125 = value__15[31:21] ^ value__15[10:0] ^ value__15[27:17];
  assign s_0__124 = value__15[20:7] ^ value__15[31:18] ^ value__15[16:3];
  assign s_1__127 = value__54[16:7] ^ value__54[18:9];
  assign s_1__126 = value__54[6:0] ^ value__54[8:2] ^ value__54[31:25];
  assign s_1__125 = value__54[31:30] ^ value__54[1:0] ^ value__54[24:23];
  assign s_1__124 = value__54[29:17] ^ value__54[31:19] ^ value__54[22:10];
  assign S1__203 = e__35[5:0] ^ e__35[10:5] ^ e__35[24:19];
  assign S1__202 = e__35[31:27] ^ e__35[4:0] ^ e__35[18:14];
  assign S1__201 = e__35[26:13] ^ e__35[31:18] ^ e__35[13:0];
  assign S1__200 = e__35[12:6] ^ e__35[17:11] ^ e__35[31:25];
  assign s_0__20 = {s_0__127, s_0__126, s_0__125, s_0__124};
  assign s_1__20 = {s_1__127, s_1__126, s_1__125, s_1__124};
  assign S0__187 = a__31[1:0] ^ a__31[12:11] ^ a__31[21:20];
  assign S0__186 = a__31[31:21] ^ a__31[10:0] ^ a__31[19:9];
  assign S0__185 = a__31[20:12] ^ a__31[31:23] ^ a__31[8:0];
  assign S0__184 = a__31[11:2] ^ a__31[22:13] ^ a__31[31:22];
  assign and_58980 = a__31 & a__30;
  assign S1__35 = {S1__203, S1__202, S1__201, S1__200};
  assign value__58 = value__12 + s_0__20;
  assign value__59 = value__39 + s_1__20;
  assign S0__31 = {S0__187, S0__186, S0__185, S0__184};
  assign maj__31 = and_58980 ^ a__31 & a__29 ^ and_58894;
  assign temp1__141 = e__32 + S1__35;
  assign ch__35 = e__35 & e__34 ^ ~(e__35 | ~e__33);
  assign value__60 = value__58 + value__59;
  assign s_0__131 = value__18[6:4] ^ value__18[17:15];
  assign s_0__130 = value__18[3:0] ^ value__18[14:11] ^ value__18[31:28];
  assign s_0__129 = value__18[31:21] ^ value__18[10:0] ^ value__18[27:17];
  assign s_0__128 = value__18[20:7] ^ value__18[31:18] ^ value__18[16:3];
  assign s_1__131 = value__57[16:7] ^ value__57[18:9];
  assign s_1__130 = value__57[6:0] ^ value__57[8:2] ^ value__57[31:25];
  assign s_1__129 = value__57[31:30] ^ value__57[1:0] ^ value__57[24:23];
  assign s_1__128 = value__57[29:17] ^ value__57[31:19] ^ value__57[22:10];
  assign temp2__31 = S0__31 + maj__31;
  assign temp1__142 = temp1__141 + ch__35;
  assign temp1__293 = value__60 + 32'h5338_0d13;
  assign s_0__21 = {s_0__131, s_0__130, s_0__129, s_0__128};
  assign s_1__21 = {s_1__131, s_1__130, s_1__129, s_1__128};
  assign a__32 = temp1__128 + temp2__31;
  assign temp1__144 = temp1__142 + temp1__293;
  assign value__61 = value__15 + s_0__21;
  assign value__62 = value__42 + s_1__21;
  assign e__36 = a__32 + temp1__144;
  assign value__63 = value__61 + value__62;
  assign S0__191 = a__32[1:0] ^ a__32[12:11] ^ a__32[21:20];
  assign S0__190 = a__32[31:21] ^ a__32[10:0] ^ a__32[19:9];
  assign S0__189 = a__32[20:12] ^ a__32[31:23] ^ a__32[8:0];
  assign S0__188 = a__32[11:2] ^ a__32[22:13] ^ a__32[31:22];
  assign and_59064 = a__32 & a__31;
  assign S1__207 = e__36[5:0] ^ e__36[10:5] ^ e__36[24:19];
  assign S1__206 = e__36[31:27] ^ e__36[4:0] ^ e__36[18:14];
  assign S1__205 = e__36[26:13] ^ e__36[31:18] ^ e__36[13:0];
  assign S1__204 = e__36[12:6] ^ e__36[17:11] ^ e__36[31:25];
  assign add_59072 = value__63[31:2] + 30'h1942_9cd5;
  assign S0__32 = {S0__191, S0__190, S0__189, S0__188};
  assign maj__32 = and_59064 ^ a__32 & a__30 ^ and_58980;
  assign S1__36 = {S1__207, S1__206, S1__205, S1__204};
  assign ch__36 = e__36 & e__35 ^ ~(e__36 | ~e__34);
  assign temp1__294 = {add_59072, value__63[1:0]};
  assign temp2__32 = S0__32 + maj__32;
  assign temp1__389 = e__33 + S1__36;
  assign temp1__390 = ch__36 + temp1__294;
  assign a__33 = temp1__132 + temp2__32;
  assign temp1__391 = temp1__389 + temp1__390;
  assign e__37 = a__33 + temp1__391;
  assign s_0__135 = value__21[6:4] ^ value__21[17:15];
  assign s_0__134 = value__21[3:0] ^ value__21[14:11] ^ value__21[31:28];
  assign s_0__133 = value__21[31:21] ^ value__21[10:0] ^ value__21[27:17];
  assign s_0__132 = value__21[20:7] ^ value__21[31:18] ^ value__21[16:3];
  assign s_1__135 = value__60[16:7] ^ value__60[18:9];
  assign s_1__134 = value__60[6:0] ^ value__60[8:2] ^ value__60[31:25];
  assign s_1__133 = value__60[31:30] ^ value__60[1:0] ^ value__60[24:23];
  assign s_1__132 = value__60[29:17] ^ value__60[31:19] ^ value__60[22:10];
  assign S1__211 = e__37[5:0] ^ e__37[10:5] ^ e__37[24:19];
  assign S1__210 = e__37[31:27] ^ e__37[4:0] ^ e__37[18:14];
  assign S1__209 = e__37[26:13] ^ e__37[31:18] ^ e__37[13:0];
  assign S1__208 = e__37[12:6] ^ e__37[17:11] ^ e__37[31:25];
  assign s_0__22 = {s_0__135, s_0__134, s_0__133, s_0__132};
  assign s_1__22 = {s_1__135, s_1__134, s_1__133, s_1__132};
  assign S0__195 = a__33[1:0] ^ a__33[12:11] ^ a__33[21:20];
  assign S0__194 = a__33[31:21] ^ a__33[10:0] ^ a__33[19:9];
  assign S0__193 = a__33[20:12] ^ a__33[31:23] ^ a__33[8:0];
  assign S0__192 = a__33[11:2] ^ a__33[22:13] ^ a__33[31:22];
  assign and_59150 = a__33 & a__32;
  assign S1__37 = {S1__211, S1__210, S1__209, S1__208};
  assign value__64 = value__18 + s_0__22;
  assign value__65 = value__45 + s_1__22;
  assign S0__33 = {S0__195, S0__194, S0__193, S0__192};
  assign maj__33 = and_59150 ^ a__33 & a__31 ^ and_59064;
  assign temp1__149 = e__34 + S1__37;
  assign ch__37 = e__37 & e__36 ^ ~(e__37 | ~e__35);
  assign value__66 = value__64 + value__65;
  assign s_0__139 = value__24[6:4] ^ value__24[17:15];
  assign s_0__138 = value__24[3:0] ^ value__24[14:11] ^ value__24[31:28];
  assign s_0__137 = value__24[31:21] ^ value__24[10:0] ^ value__24[27:17];
  assign s_0__136 = value__24[20:7] ^ value__24[31:18] ^ value__24[16:3];
  assign s_1__139 = value__63[16:7] ^ value__63[18:9];
  assign s_1__138 = value__63[6:0] ^ value__63[8:2] ^ value__63[31:25];
  assign s_1__137 = value__63[31:30] ^ value__63[1:0] ^ value__63[24:23];
  assign s_1__136 = value__63[29:17] ^ value__63[31:19] ^ value__63[22:10];
  assign temp2__33 = S0__33 + maj__33;
  assign temp1__150 = temp1__149 + ch__37;
  assign temp1__295 = value__66 + 32'h766a_0abb;
  assign s_0__23 = {s_0__139, s_0__138, s_0__137, s_0__136};
  assign s_1__23 = {s_1__139, s_1__138, s_1__137, s_1__136};
  assign a__34 = temp1__397 + temp2__33;
  assign temp1__152 = temp1__150 + temp1__295;
  assign value__67 = value__21 + s_0__23;
  assign value__68 = value__48 + s_1__23;
  assign e__38 = a__34 + temp1__152;
  assign value__69 = value__67 + value__68;
  assign S0__199 = a__34[1:0] ^ a__34[12:11] ^ a__34[21:20];
  assign S0__198 = a__34[31:21] ^ a__34[10:0] ^ a__34[19:9];
  assign S0__197 = a__34[20:12] ^ a__34[31:23] ^ a__34[8:0];
  assign S0__196 = a__34[11:2] ^ a__34[22:13] ^ a__34[31:22];
  assign and_59234 = a__34 & a__33;
  assign S1__215 = e__38[5:0] ^ e__38[10:5] ^ e__38[24:19];
  assign S1__214 = e__38[31:27] ^ e__38[4:0] ^ e__38[18:14];
  assign S1__213 = e__38[26:13] ^ e__38[31:18] ^ e__38[13:0];
  assign S1__212 = e__38[12:6] ^ e__38[17:11] ^ e__38[31:25];
  assign add_59242 = value__69[31:1] + 31'h40e1_6497;
  assign S0__34 = {S0__199, S0__198, S0__197, S0__196};
  assign maj__34 = and_59234 ^ a__34 & a__32 ^ and_59150;
  assign S1__38 = {S1__215, S1__214, S1__213, S1__212};
  assign ch__38 = e__38 & e__37 ^ ~(e__38 | ~e__36);
  assign temp1__296 = {add_59242, value__69[0]};
  assign temp2__34 = S0__34 + maj__34;
  assign temp1__386 = e__35 + S1__38;
  assign temp1__387 = ch__38 + temp1__296;
  assign a__35 = temp1__394 + temp2__34;
  assign temp1__388 = temp1__386 + temp1__387;
  assign e__39 = a__35 + temp1__388;
  assign s_0__143 = value__27[6:4] ^ value__27[17:15];
  assign s_0__142 = value__27[3:0] ^ value__27[14:11] ^ value__27[31:28];
  assign s_0__141 = value__27[31:21] ^ value__27[10:0] ^ value__27[27:17];
  assign s_0__140 = value__27[20:7] ^ value__27[31:18] ^ value__27[16:3];
  assign s_1__143 = value__66[16:7] ^ value__66[18:9];
  assign s_1__142 = value__66[6:0] ^ value__66[8:2] ^ value__66[31:25];
  assign s_1__141 = value__66[31:30] ^ value__66[1:0] ^ value__66[24:23];
  assign s_1__140 = value__66[29:17] ^ value__66[31:19] ^ value__66[22:10];
  assign S1__219 = e__39[5:0] ^ e__39[10:5] ^ e__39[24:19];
  assign S1__218 = e__39[31:27] ^ e__39[4:0] ^ e__39[18:14];
  assign S1__217 = e__39[26:13] ^ e__39[31:18] ^ e__39[13:0];
  assign S1__216 = e__39[12:6] ^ e__39[17:11] ^ e__39[31:25];
  assign s_0__24 = {s_0__143, s_0__142, s_0__141, s_0__140};
  assign s_1__24 = {s_1__143, s_1__142, s_1__141, s_1__140};
  assign S0__203 = a__35[1:0] ^ a__35[12:11] ^ a__35[21:20];
  assign S0__202 = a__35[31:21] ^ a__35[10:0] ^ a__35[19:9];
  assign S0__201 = a__35[20:12] ^ a__35[31:23] ^ a__35[8:0];
  assign S0__200 = a__35[11:2] ^ a__35[22:13] ^ a__35[31:22];
  assign and_59320 = a__35 & a__34;
  assign S1__39 = {S1__219, S1__218, S1__217, S1__216};
  assign value__70 = value__24 + s_0__24;
  assign value__71 = value__51 + s_1__24;
  assign S0__35 = {S0__203, S0__202, S0__201, S0__200};
  assign maj__35 = and_59320 ^ a__35 & a__33 ^ and_59234;
  assign temp1__157 = e__36 + S1__39;
  assign ch__39 = e__39 & e__38 ^ ~(e__39 | ~e__37);
  assign value__72 = value__70 + value__71;
  assign temp2__35 = S0__35 + maj__35;
  assign temp1__158 = temp1__157 + ch__39;
  assign temp1__297 = value__72 + 32'h9272_2c85;
  assign a__36 = temp1__144 + temp2__35;
  assign temp1__160 = temp1__158 + temp1__297;
  assign e__40 = a__36 + temp1__160;
  assign s_0__147 = value__30[6:4] ^ value__30[17:15];
  assign s_0__146 = value__30[3:0] ^ value__30[14:11] ^ value__30[31:28];
  assign s_0__145 = value__30[31:21] ^ value__30[10:0] ^ value__30[27:17];
  assign s_0__144 = value__30[20:7] ^ value__30[31:18] ^ value__30[16:3];
  assign s_1__147 = value__69[16:7] ^ value__69[18:9];
  assign s_1__146 = value__69[6:0] ^ value__69[8:2] ^ value__69[31:25];
  assign s_1__145 = value__69[31:30] ^ value__69[1:0] ^ value__69[24:23];
  assign s_1__144 = value__69[29:17] ^ value__69[31:19] ^ value__69[22:10];
  assign S1__223 = e__40[5:0] ^ e__40[10:5] ^ e__40[24:19];
  assign S1__222 = e__40[31:27] ^ e__40[4:0] ^ e__40[18:14];
  assign S1__221 = e__40[26:13] ^ e__40[31:18] ^ e__40[13:0];
  assign S1__220 = e__40[12:6] ^ e__40[17:11] ^ e__40[31:25];
  assign s_0__25 = {s_0__147, s_0__146, s_0__145, s_0__144};
  assign s_1__25 = {s_1__147, s_1__146, s_1__145, s_1__144};
  assign S0__207 = a__36[1:0] ^ a__36[12:11] ^ a__36[21:20];
  assign S0__206 = a__36[31:21] ^ a__36[10:0] ^ a__36[19:9];
  assign S0__205 = a__36[20:12] ^ a__36[31:23] ^ a__36[8:0];
  assign S0__204 = a__36[11:2] ^ a__36[22:13] ^ a__36[31:22];
  assign and_59404 = a__36 & a__35;
  assign S1__40 = {S1__223, S1__222, S1__221, S1__220};
  assign value__73 = value__27 + s_0__25;
  assign value__74 = value__54 + s_1__25;
  assign S0__36 = {S0__207, S0__206, S0__205, S0__204};
  assign maj__36 = and_59404 ^ a__36 & a__34 ^ and_59320;
  assign temp1__161 = e__37 + S1__40;
  assign ch__40 = e__40 & e__39 ^ ~(e__40 | ~e__38);
  assign value__75 = value__73 + value__74;
  assign temp2__36 = S0__36 + maj__36;
  assign temp1__162 = temp1__161 + ch__40;
  assign temp1__298 = value__75 + 32'ha2bf_e8a1;
  assign a__37 = temp1__391 + temp2__36;
  assign temp1__164 = temp1__162 + temp1__298;
  assign e__41 = a__37 + temp1__164;
  assign s_0__151 = value__33[6:4] ^ value__33[17:15];
  assign s_0__150 = value__33[3:0] ^ value__33[14:11] ^ value__33[31:28];
  assign s_0__149 = value__33[31:21] ^ value__33[10:0] ^ value__33[27:17];
  assign s_0__148 = value__33[20:7] ^ value__33[31:18] ^ value__33[16:3];
  assign s_1__151 = value__72[16:7] ^ value__72[18:9];
  assign s_1__150 = value__72[6:0] ^ value__72[8:2] ^ value__72[31:25];
  assign s_1__149 = value__72[31:30] ^ value__72[1:0] ^ value__72[24:23];
  assign s_1__148 = value__72[29:17] ^ value__72[31:19] ^ value__72[22:10];
  assign S1__227 = e__41[5:0] ^ e__41[10:5] ^ e__41[24:19];
  assign S1__226 = e__41[31:27] ^ e__41[4:0] ^ e__41[18:14];
  assign S1__225 = e__41[26:13] ^ e__41[31:18] ^ e__41[13:0];
  assign S1__224 = e__41[12:6] ^ e__41[17:11] ^ e__41[31:25];
  assign s_0__26 = {s_0__151, s_0__150, s_0__149, s_0__148};
  assign s_1__26 = {s_1__151, s_1__150, s_1__149, s_1__148};
  assign S0__211 = a__37[1:0] ^ a__37[12:11] ^ a__37[21:20];
  assign S0__210 = a__37[31:21] ^ a__37[10:0] ^ a__37[19:9];
  assign S0__209 = a__37[20:12] ^ a__37[31:23] ^ a__37[8:0];
  assign S0__208 = a__37[11:2] ^ a__37[22:13] ^ a__37[31:22];
  assign and_59488 = a__37 & a__36;
  assign S1__41 = {S1__227, S1__226, S1__225, S1__224};
  assign value__76 = value__30 + s_0__26;
  assign value__77 = value__57 + s_1__26;
  assign S0__37 = {S0__211, S0__210, S0__209, S0__208};
  assign maj__37 = and_59488 ^ a__37 & a__35 ^ and_59404;
  assign temp1__165 = e__38 + S1__41;
  assign ch__41 = e__41 & e__40 ^ ~(e__41 | ~e__39);
  assign value__78 = value__76 + value__77;
  assign s_0__155 = value__36[6:4] ^ value__36[17:15];
  assign s_0__154 = value__36[3:0] ^ value__36[14:11] ^ value__36[31:28];
  assign s_0__153 = value__36[31:21] ^ value__36[10:0] ^ value__36[27:17];
  assign s_0__152 = value__36[20:7] ^ value__36[31:18] ^ value__36[16:3];
  assign s_1__155 = value__75[16:7] ^ value__75[18:9];
  assign s_1__154 = value__75[6:0] ^ value__75[8:2] ^ value__75[31:25];
  assign s_1__153 = value__75[31:30] ^ value__75[1:0] ^ value__75[24:23];
  assign s_1__152 = value__75[29:17] ^ value__75[31:19] ^ value__75[22:10];
  assign temp2__37 = S0__37 + maj__37;
  assign temp1__166 = temp1__165 + ch__41;
  assign temp1__299 = value__78 + 32'ha81a_664b;
  assign s_0__27 = {s_0__155, s_0__154, s_0__153, s_0__152};
  assign s_1__27 = {s_1__155, s_1__154, s_1__153, s_1__152};
  assign a__38 = temp1__152 + temp2__37;
  assign temp1__168 = temp1__166 + temp1__299;
  assign value__79 = value__33 + s_0__27;
  assign value__80 = value__60 + s_1__27;
  assign e__42 = a__38 + temp1__168;
  assign value__81 = value__79 + value__80;
  assign S0__215 = a__38[1:0] ^ a__38[12:11] ^ a__38[21:20];
  assign S0__214 = a__38[31:21] ^ a__38[10:0] ^ a__38[19:9];
  assign S0__213 = a__38[20:12] ^ a__38[31:23] ^ a__38[8:0];
  assign S0__212 = a__38[11:2] ^ a__38[22:13] ^ a__38[31:22];
  assign and_59573 = a__38 & a__37;
  assign S1__231 = e__42[5:0] ^ e__42[10:5] ^ e__42[24:19];
  assign S1__230 = e__42[31:27] ^ e__42[4:0] ^ e__42[18:14];
  assign S1__229 = e__42[26:13] ^ e__42[31:18] ^ e__42[13:0];
  assign S1__228 = e__42[12:6] ^ e__42[17:11] ^ e__42[31:25];
  assign add_59581 = value__81[31:4] + 28'hc24_b8b7;
  assign S0__38 = {S0__215, S0__214, S0__213, S0__212};
  assign maj__38 = and_59573 ^ a__38 & a__36 ^ and_59488;
  assign S1__42 = {S1__231, S1__230, S1__229, S1__228};
  assign ch__42 = e__42 & e__41 ^ ~(e__42 | ~e__40);
  assign temp1__300 = {add_59581, value__81[3:0]};
  assign temp2__38 = S0__38 + maj__38;
  assign temp1__383 = e__39 + S1__42;
  assign temp1__384 = ch__42 + temp1__300;
  assign a__39 = temp1__388 + temp2__38;
  assign temp1__385 = temp1__383 + temp1__384;
  assign e__43 = a__39 + temp1__385;
  assign s_0__159 = value__39[6:4] ^ value__39[17:15];
  assign s_0__158 = value__39[3:0] ^ value__39[14:11] ^ value__39[31:28];
  assign s_0__157 = value__39[31:21] ^ value__39[10:0] ^ value__39[27:17];
  assign s_0__156 = value__39[20:7] ^ value__39[31:18] ^ value__39[16:3];
  assign s_1__159 = value__78[16:7] ^ value__78[18:9];
  assign s_1__158 = value__78[6:0] ^ value__78[8:2] ^ value__78[31:25];
  assign s_1__157 = value__78[31:30] ^ value__78[1:0] ^ value__78[24:23];
  assign s_1__156 = value__78[29:17] ^ value__78[31:19] ^ value__78[22:10];
  assign S1__235 = e__43[5:0] ^ e__43[10:5] ^ e__43[24:19];
  assign S1__234 = e__43[31:27] ^ e__43[4:0] ^ e__43[18:14];
  assign S1__233 = e__43[26:13] ^ e__43[31:18] ^ e__43[13:0];
  assign S1__232 = e__43[12:6] ^ e__43[17:11] ^ e__43[31:25];
  assign s_0__28 = {s_0__159, s_0__158, s_0__157, s_0__156};
  assign s_1__28 = {s_1__159, s_1__158, s_1__157, s_1__156};
  assign S0__219 = a__39[1:0] ^ a__39[12:11] ^ a__39[21:20];
  assign S0__218 = a__39[31:21] ^ a__39[10:0] ^ a__39[19:9];
  assign S0__217 = a__39[20:12] ^ a__39[31:23] ^ a__39[8:0];
  assign S0__216 = a__39[11:2] ^ a__39[22:13] ^ a__39[31:22];
  assign and_59659 = a__39 & a__38;
  assign S1__43 = {S1__235, S1__234, S1__233, S1__232};
  assign value__82 = value__36 + s_0__28;
  assign value__83 = value__63 + s_1__28;
  assign S0__39 = {S0__219, S0__218, S0__217, S0__216};
  assign maj__39 = and_59659 ^ a__39 & a__37 ^ and_59573;
  assign temp1__173 = e__40 + S1__43;
  assign ch__43 = e__43 & e__42 ^ ~(e__43 | ~e__41);
  assign value__84 = value__82 + value__83;
  assign temp2__39 = S0__39 + maj__39;
  assign temp1__174 = temp1__173 + ch__43;
  assign temp1__301 = value__84 + 32'hc76c_51a3;
  assign a__40 = temp1__160 + temp2__39;
  assign temp1__176 = temp1__174 + temp1__301;
  assign e__44 = a__40 + temp1__176;
  assign s_0__163 = value__42[6:4] ^ value__42[17:15];
  assign s_0__162 = value__42[3:0] ^ value__42[14:11] ^ value__42[31:28];
  assign s_0__161 = value__42[31:21] ^ value__42[10:0] ^ value__42[27:17];
  assign s_0__160 = value__42[20:7] ^ value__42[31:18] ^ value__42[16:3];
  assign s_1__163 = value__81[16:7] ^ value__81[18:9];
  assign s_1__162 = value__81[6:0] ^ value__81[8:2] ^ value__81[31:25];
  assign s_1__161 = value__81[31:30] ^ value__81[1:0] ^ value__81[24:23];
  assign s_1__160 = value__81[29:17] ^ value__81[31:19] ^ value__81[22:10];
  assign S1__239 = e__44[5:0] ^ e__44[10:5] ^ e__44[24:19];
  assign S1__238 = e__44[31:27] ^ e__44[4:0] ^ e__44[18:14];
  assign S1__237 = e__44[26:13] ^ e__44[31:18] ^ e__44[13:0];
  assign S1__236 = e__44[12:6] ^ e__44[17:11] ^ e__44[31:25];
  assign s_0__29 = {s_0__163, s_0__162, s_0__161, s_0__160};
  assign s_1__29 = {s_1__163, s_1__162, s_1__161, s_1__160};
  assign S0__223 = a__40[1:0] ^ a__40[12:11] ^ a__40[21:20];
  assign S0__222 = a__40[31:21] ^ a__40[10:0] ^ a__40[19:9];
  assign S0__221 = a__40[20:12] ^ a__40[31:23] ^ a__40[8:0];
  assign S0__220 = a__40[11:2] ^ a__40[22:13] ^ a__40[31:22];
  assign and_59743 = a__40 & a__39;
  assign S1__44 = {S1__239, S1__238, S1__237, S1__236};
  assign value__85 = value__39 + s_0__29;
  assign value__86 = value__66 + s_1__29;
  assign S0__40 = {S0__223, S0__222, S0__221, S0__220};
  assign maj__40 = and_59743 ^ a__40 & a__38 ^ and_59659;
  assign temp1__177 = e__41 + S1__44;
  assign ch__44 = e__44 & e__43 ^ ~(e__44 | ~e__42);
  assign value__87 = value__85 + value__86;
  assign s_0__167 = value__45[6:4] ^ value__45[17:15];
  assign s_0__166 = value__45[3:0] ^ value__45[14:11] ^ value__45[31:28];
  assign s_0__165 = value__45[31:21] ^ value__45[10:0] ^ value__45[27:17];
  assign s_0__164 = value__45[20:7] ^ value__45[31:18] ^ value__45[16:3];
  assign s_1__167 = value__84[16:7] ^ value__84[18:9];
  assign s_1__166 = value__84[6:0] ^ value__84[8:2] ^ value__84[31:25];
  assign s_1__165 = value__84[31:30] ^ value__84[1:0] ^ value__84[24:23];
  assign s_1__164 = value__84[29:17] ^ value__84[31:19] ^ value__84[22:10];
  assign temp2__40 = S0__40 + maj__40;
  assign temp1__178 = temp1__177 + ch__44;
  assign temp1__302 = value__87 + 32'hd192_e819;
  assign s_0__30 = {s_0__167, s_0__166, s_0__165, s_0__164};
  assign s_1__30 = {s_1__167, s_1__166, s_1__165, s_1__164};
  assign a__41 = temp1__164 + temp2__40;
  assign temp1__180 = temp1__178 + temp1__302;
  assign value__88 = value__42 + s_0__30;
  assign value__89 = value__69 + s_1__30;
  assign e__45 = a__41 + temp1__180;
  assign value__90 = value__88 + value__89;
  assign S0__227 = a__41[1:0] ^ a__41[12:11] ^ a__41[21:20];
  assign S0__226 = a__41[31:21] ^ a__41[10:0] ^ a__41[19:9];
  assign S0__225 = a__41[20:12] ^ a__41[31:23] ^ a__41[8:0];
  assign S0__224 = a__41[11:2] ^ a__41[22:13] ^ a__41[31:22];
  assign and_59828 = a__41 & a__40;
  assign S1__243 = e__45[5:0] ^ e__45[10:5] ^ e__45[24:19];
  assign S1__242 = e__45[31:27] ^ e__45[4:0] ^ e__45[18:14];
  assign S1__241 = e__45[26:13] ^ e__45[31:18] ^ e__45[13:0];
  assign S1__240 = e__45[12:6] ^ e__45[17:11] ^ e__45[31:25];
  assign add_59836 = value__90[31:2] + 30'h35a6_4189;
  assign S0__41 = {S0__227, S0__226, S0__225, S0__224};
  assign maj__41 = and_59828 ^ a__41 & a__39 ^ and_59743;
  assign S1__45 = {S1__243, S1__242, S1__241, S1__240};
  assign ch__45 = e__45 & e__44 ^ ~(e__45 | ~e__43);
  assign temp1__303 = {add_59836, value__90[1:0]};
  assign temp2__41 = S0__41 + maj__41;
  assign temp1__380 = e__42 + S1__45;
  assign temp1__381 = ch__45 + temp1__303;
  assign a__42 = temp1__168 + temp2__41;
  assign temp1__382 = temp1__380 + temp1__381;
  assign e__46 = a__42 + temp1__382;
  assign s_0__171 = value__48[6:4] ^ value__48[17:15];
  assign s_0__170 = value__48[3:0] ^ value__48[14:11] ^ value__48[31:28];
  assign s_0__169 = value__48[31:21] ^ value__48[10:0] ^ value__48[27:17];
  assign s_0__168 = value__48[20:7] ^ value__48[31:18] ^ value__48[16:3];
  assign s_1__171 = value__87[16:7] ^ value__87[18:9];
  assign s_1__170 = value__87[6:0] ^ value__87[8:2] ^ value__87[31:25];
  assign s_1__169 = value__87[31:30] ^ value__87[1:0] ^ value__87[24:23];
  assign s_1__168 = value__87[29:17] ^ value__87[31:19] ^ value__87[22:10];
  assign S1__247 = e__46[5:0] ^ e__46[10:5] ^ e__46[24:19];
  assign S1__246 = e__46[31:27] ^ e__46[4:0] ^ e__46[18:14];
  assign S1__245 = e__46[26:13] ^ e__46[31:18] ^ e__46[13:0];
  assign S1__244 = e__46[12:6] ^ e__46[17:11] ^ e__46[31:25];
  assign s_0__31 = {s_0__171, s_0__170, s_0__169, s_0__168};
  assign s_1__31 = {s_1__171, s_1__170, s_1__169, s_1__168};
  assign S0__231 = a__42[1:0] ^ a__42[12:11] ^ a__42[21:20];
  assign S0__230 = a__42[31:21] ^ a__42[10:0] ^ a__42[19:9];
  assign S0__229 = a__42[20:12] ^ a__42[31:23] ^ a__42[8:0];
  assign S0__228 = a__42[11:2] ^ a__42[22:13] ^ a__42[31:22];
  assign and_59914 = a__42 & a__41;
  assign S1__46 = {S1__247, S1__246, S1__245, S1__244};
  assign value__91 = value__45 + s_0__31;
  assign value__92 = value__72 + s_1__31;
  assign S0__42 = {S0__231, S0__230, S0__229, S0__228};
  assign maj__42 = and_59914 ^ a__42 & a__40 ^ and_59828;
  assign temp1__185 = e__43 + S1__46;
  assign ch__46 = e__46 & e__45 ^ ~(e__46 | ~e__44);
  assign value__93 = value__91 + value__92;
  assign s_0__175 = value__51[6:4] ^ value__51[17:15];
  assign s_0__174 = value__51[3:0] ^ value__51[14:11] ^ value__51[31:28];
  assign s_0__173 = value__51[31:21] ^ value__51[10:0] ^ value__51[27:17];
  assign s_0__172 = value__51[20:7] ^ value__51[31:18] ^ value__51[16:3];
  assign s_1__175 = value__90[16:7] ^ value__90[18:9];
  assign s_1__174 = value__90[6:0] ^ value__90[8:2] ^ value__90[31:25];
  assign s_1__173 = value__90[31:30] ^ value__90[1:0] ^ value__90[24:23];
  assign s_1__172 = value__90[29:17] ^ value__90[31:19] ^ value__90[22:10];
  assign temp2__42 = S0__42 + maj__42;
  assign temp1__186 = temp1__185 + ch__46;
  assign temp1__304 = value__93 + 32'hf40e_3585;
  assign s_0__32 = {s_0__175, s_0__174, s_0__173, s_0__172};
  assign s_1__32 = {s_1__175, s_1__174, s_1__173, s_1__172};
  assign a__43 = temp1__385 + temp2__42;
  assign temp1__188 = temp1__186 + temp1__304;
  assign value__94 = value__48 + s_0__32;
  assign value__95 = value__75 + s_1__32;
  assign e__47 = a__43 + temp1__188;
  assign value__96 = value__94 + value__95;
  assign S0__235 = a__43[1:0] ^ a__43[12:11] ^ a__43[21:20];
  assign S0__234 = a__43[31:21] ^ a__43[10:0] ^ a__43[19:9];
  assign S0__233 = a__43[20:12] ^ a__43[31:23] ^ a__43[8:0];
  assign S0__232 = a__43[11:2] ^ a__43[22:13] ^ a__43[31:22];
  assign and_59998 = a__43 & a__42;
  assign S1__251 = e__47[5:0] ^ e__47[10:5] ^ e__47[24:19];
  assign S1__250 = e__47[31:27] ^ e__47[4:0] ^ e__47[18:14];
  assign S1__249 = e__47[26:13] ^ e__47[31:18] ^ e__47[13:0];
  assign S1__248 = e__47[12:6] ^ e__47[17:11] ^ e__47[31:25];
  assign add_60006 = value__96[31:4] + 28'h106_aa07;
  assign S0__43 = {S0__235, S0__234, S0__233, S0__232};
  assign maj__43 = and_59998 ^ a__43 & a__41 ^ and_59914;
  assign S1__47 = {S1__251, S1__250, S1__249, S1__248};
  assign ch__47 = e__47 & e__46 ^ ~(e__47 | ~e__45);
  assign temp1__305 = {add_60006, value__96[3:0]};
  assign s_0__179 = value__54[6:4] ^ value__54[17:15];
  assign s_0__178 = value__54[3:0] ^ value__54[14:11] ^ value__54[31:28];
  assign s_0__177 = value__54[31:21] ^ value__54[10:0] ^ value__54[27:17];
  assign s_0__176 = value__54[20:7] ^ value__54[31:18] ^ value__54[16:3];
  assign s_1__179 = value__93[16:7] ^ value__93[18:9];
  assign s_1__178 = value__93[6:0] ^ value__93[8:2] ^ value__93[31:25];
  assign s_1__177 = value__93[31:30] ^ value__93[1:0] ^ value__93[24:23];
  assign s_1__176 = value__93[29:17] ^ value__93[31:19] ^ value__93[22:10];
  assign temp2__43 = S0__43 + maj__43;
  assign temp1__377 = e__44 + S1__47;
  assign temp1__378 = ch__47 + temp1__305;
  assign s_0__33 = {s_0__179, s_0__178, s_0__177, s_0__176};
  assign s_1__33 = {s_1__179, s_1__178, s_1__177, s_1__176};
  assign a__44 = temp1__176 + temp2__43;
  assign temp1__379 = temp1__377 + temp1__378;
  assign value__97 = value__51 + s_0__33;
  assign value__98 = value__78 + s_1__33;
  assign e__48 = a__44 + temp1__379;
  assign value__99 = value__97 + value__98;
  assign S0__239 = a__44[1:0] ^ a__44[12:11] ^ a__44[21:20];
  assign S0__238 = a__44[31:21] ^ a__44[10:0] ^ a__44[19:9];
  assign S0__237 = a__44[20:12] ^ a__44[31:23] ^ a__44[8:0];
  assign S0__236 = a__44[11:2] ^ a__44[22:13] ^ a__44[31:22];
  assign and_60085 = a__44 & a__43;
  assign S1__255 = e__48[5:0] ^ e__48[10:5] ^ e__48[24:19];
  assign S1__254 = e__48[31:27] ^ e__48[4:0] ^ e__48[18:14];
  assign S1__253 = e__48[26:13] ^ e__48[31:18] ^ e__48[13:0];
  assign S1__252 = e__48[12:6] ^ e__48[17:11] ^ e__48[31:25];
  assign add_60093 = value__99[31:1] + 31'h0cd2_608b;
  assign S0__44 = {S0__239, S0__238, S0__237, S0__236};
  assign maj__44 = and_60085 ^ a__44 & a__42 ^ and_59998;
  assign S1__48 = {S1__255, S1__254, S1__253, S1__252};
  assign ch__48 = e__48 & e__47 ^ ~(e__48 | ~e__46);
  assign temp1__306 = {add_60093, value__99[0]};
  assign s_0__183 = value__57[6:4] ^ value__57[17:15];
  assign s_0__182 = value__57[3:0] ^ value__57[14:11] ^ value__57[31:28];
  assign s_0__181 = value__57[31:21] ^ value__57[10:0] ^ value__57[27:17];
  assign s_0__180 = value__57[20:7] ^ value__57[31:18] ^ value__57[16:3];
  assign s_1__183 = value__96[16:7] ^ value__96[18:9];
  assign s_1__182 = value__96[6:0] ^ value__96[8:2] ^ value__96[31:25];
  assign s_1__181 = value__96[31:30] ^ value__96[1:0] ^ value__96[24:23];
  assign s_1__180 = value__96[29:17] ^ value__96[31:19] ^ value__96[22:10];
  assign temp2__44 = S0__44 + maj__44;
  assign temp1__374 = e__45 + S1__48;
  assign temp1__375 = ch__48 + temp1__306;
  assign s_0__34 = {s_0__183, s_0__182, s_0__181, s_0__180};
  assign s_1__34 = {s_1__183, s_1__182, s_1__181, s_1__180};
  assign a__45 = temp1__180 + temp2__44;
  assign temp1__376 = temp1__374 + temp1__375;
  assign value__100 = value__54 + s_0__34;
  assign value__101 = value__81 + s_1__34;
  assign e__49 = a__45 + temp1__376;
  assign value__102 = value__100 + value__101;
  assign S0__243 = a__45[1:0] ^ a__45[12:11] ^ a__45[21:20];
  assign S0__242 = a__45[31:21] ^ a__45[10:0] ^ a__45[19:9];
  assign S0__241 = a__45[20:12] ^ a__45[31:23] ^ a__45[8:0];
  assign S0__240 = a__45[11:2] ^ a__45[22:13] ^ a__45[31:22];
  assign and_60172 = a__45 & a__44;
  assign S1__259 = e__49[5:0] ^ e__49[10:5] ^ e__49[24:19];
  assign S1__258 = e__49[31:27] ^ e__49[4:0] ^ e__49[18:14];
  assign S1__257 = e__49[26:13] ^ e__49[31:18] ^ e__49[13:0];
  assign S1__256 = e__49[12:6] ^ e__49[17:11] ^ e__49[31:25];
  assign add_60180 = value__102[31:3] + 29'h03c6_ed81;
  assign S0__45 = {S0__243, S0__242, S0__241, S0__240};
  assign maj__45 = and_60172 ^ a__45 & a__43 ^ and_60085;
  assign S1__49 = {S1__259, S1__258, S1__257, S1__256};
  assign ch__49 = e__49 & e__48 ^ ~(e__49 | ~e__47);
  assign temp1__307 = {add_60180, value__102[2:0]};
  assign s_0__187 = value__60[6:4] ^ value__60[17:15];
  assign s_0__186 = value__60[3:0] ^ value__60[14:11] ^ value__60[31:28];
  assign s_0__185 = value__60[31:21] ^ value__60[10:0] ^ value__60[27:17];
  assign s_0__184 = value__60[20:7] ^ value__60[31:18] ^ value__60[16:3];
  assign s_1__187 = value__99[16:7] ^ value__99[18:9];
  assign s_1__186 = value__99[6:0] ^ value__99[8:2] ^ value__99[31:25];
  assign s_1__185 = value__99[31:30] ^ value__99[1:0] ^ value__99[24:23];
  assign s_1__184 = value__99[29:17] ^ value__99[31:19] ^ value__99[22:10];
  assign temp2__45 = S0__45 + maj__45;
  assign temp1__371 = e__46 + S1__49;
  assign temp1__372 = ch__49 + temp1__307;
  assign s_0__35 = {s_0__187, s_0__186, s_0__185, s_0__184};
  assign s_1__35 = {s_1__187, s_1__186, s_1__185, s_1__184};
  assign a__46 = temp1__382 + temp2__45;
  assign temp1__373 = temp1__371 + temp1__372;
  assign value__103 = value__57 + s_0__35;
  assign value__104 = value__84 + s_1__35;
  assign e__50 = a__46 + temp1__373;
  assign value__105 = value__103 + value__104;
  assign S0__247 = a__46[1:0] ^ a__46[12:11] ^ a__46[21:20];
  assign S0__246 = a__46[31:21] ^ a__46[10:0] ^ a__46[19:9];
  assign S0__245 = a__46[20:12] ^ a__46[31:23] ^ a__46[8:0];
  assign S0__244 = a__46[11:2] ^ a__46[22:13] ^ a__46[31:22];
  assign and_60259 = a__46 & a__45;
  assign S1__263 = e__50[5:0] ^ e__50[10:5] ^ e__50[24:19];
  assign S1__262 = e__50[31:27] ^ e__50[4:0] ^ e__50[18:14];
  assign S1__261 = e__50[26:13] ^ e__50[31:18] ^ e__50[13:0];
  assign S1__260 = e__50[12:6] ^ e__50[17:11] ^ e__50[31:25];
  assign add_60267 = value__105[31:2] + 30'h09d2_1dd3;
  assign S0__46 = {S0__247, S0__246, S0__245, S0__244};
  assign maj__46 = and_60259 ^ a__46 & a__44 ^ and_60172;
  assign S1__50 = {S1__263, S1__262, S1__261, S1__260};
  assign ch__50 = e__50 & e__49 ^ ~(e__50 | ~e__48);
  assign temp1__308 = {add_60267, value__105[1:0]};
  assign temp2__46 = S0__46 + maj__46;
  assign temp1__368 = e__47 + S1__50;
  assign temp1__369 = ch__50 + temp1__308;
  assign a__47 = temp1__188 + temp2__46;
  assign temp1__370 = temp1__368 + temp1__369;
  assign e__51 = a__47 + temp1__370;
  assign s_0__191 = value__63[6:4] ^ value__63[17:15];
  assign s_0__190 = value__63[3:0] ^ value__63[14:11] ^ value__63[31:28];
  assign s_0__189 = value__63[31:21] ^ value__63[10:0] ^ value__63[27:17];
  assign s_0__188 = value__63[20:7] ^ value__63[31:18] ^ value__63[16:3];
  assign s_1__191 = value__102[16:7] ^ value__102[18:9];
  assign s_1__190 = value__102[6:0] ^ value__102[8:2] ^ value__102[31:25];
  assign s_1__189 = value__102[31:30] ^ value__102[1:0] ^ value__102[24:23];
  assign s_1__188 = value__102[29:17] ^ value__102[31:19] ^ value__102[22:10];
  assign S1__267 = e__51[5:0] ^ e__51[10:5] ^ e__51[24:19];
  assign S1__266 = e__51[31:27] ^ e__51[4:0] ^ e__51[18:14];
  assign S1__265 = e__51[26:13] ^ e__51[31:18] ^ e__51[13:0];
  assign S1__264 = e__51[12:6] ^ e__51[17:11] ^ e__51[31:25];
  assign s_0__36 = {s_0__191, s_0__190, s_0__189, s_0__188};
  assign s_1__36 = {s_1__191, s_1__190, s_1__189, s_1__188};
  assign S0__251 = a__47[1:0] ^ a__47[12:11] ^ a__47[21:20];
  assign S0__250 = a__47[31:21] ^ a__47[10:0] ^ a__47[19:9];
  assign S0__249 = a__47[20:12] ^ a__47[31:23] ^ a__47[8:0];
  assign S0__248 = a__47[11:2] ^ a__47[22:13] ^ a__47[31:22];
  assign and_60345 = a__47 & a__46;
  assign S1__51 = {S1__267, S1__266, S1__265, S1__264};
  assign value__106 = value__60 + s_0__36;
  assign value__107 = value__87 + s_1__36;
  assign S0__47 = {S0__251, S0__250, S0__249, S0__248};
  assign maj__47 = and_60345 ^ a__47 & a__45 ^ and_60259;
  assign temp1__205 = e__48 + S1__51;
  assign ch__51 = e__51 & e__50 ^ ~(e__51 | ~e__49);
  assign value__108 = value__106 + value__107;
  assign temp2__47 = S0__47 + maj__47;
  assign temp1__206 = temp1__205 + ch__51;
  assign temp1__309 = value__108 + 32'h34b0_bcb5;
  assign a__48 = temp1__379 + temp2__47;
  assign temp1__208 = temp1__206 + temp1__309;
  assign e__52 = a__48 + temp1__208;
  assign s_0__195 = value__66[6:4] ^ value__66[17:15];
  assign s_0__194 = value__66[3:0] ^ value__66[14:11] ^ value__66[31:28];
  assign s_0__193 = value__66[31:21] ^ value__66[10:0] ^ value__66[27:17];
  assign s_0__192 = value__66[20:7] ^ value__66[31:18] ^ value__66[16:3];
  assign s_1__195 = value__105[16:7] ^ value__105[18:9];
  assign s_1__194 = value__105[6:0] ^ value__105[8:2] ^ value__105[31:25];
  assign s_1__193 = value__105[31:30] ^ value__105[1:0] ^ value__105[24:23];
  assign s_1__192 = value__105[29:17] ^ value__105[31:19] ^ value__105[22:10];
  assign S1__271 = e__52[5:0] ^ e__52[10:5] ^ e__52[24:19];
  assign S1__270 = e__52[31:27] ^ e__52[4:0] ^ e__52[18:14];
  assign S1__269 = e__52[26:13] ^ e__52[31:18] ^ e__52[13:0];
  assign S1__268 = e__52[12:6] ^ e__52[17:11] ^ e__52[31:25];
  assign s_0__37 = {s_0__195, s_0__194, s_0__193, s_0__192};
  assign s_1__37 = {s_1__195, s_1__194, s_1__193, s_1__192};
  assign S0__255 = a__48[1:0] ^ a__48[12:11] ^ a__48[21:20];
  assign S0__254 = a__48[31:21] ^ a__48[10:0] ^ a__48[19:9];
  assign S0__253 = a__48[20:12] ^ a__48[31:23] ^ a__48[8:0];
  assign S0__252 = a__48[11:2] ^ a__48[22:13] ^ a__48[31:22];
  assign and_60428 = a__48 & a__47;
  assign S1__52 = {S1__271, S1__270, S1__269, S1__268};
  assign value__109 = value__63 + s_0__37;
  assign value__110 = value__90 + s_1__37;
  assign S0__48 = {S0__255, S0__254, S0__253, S0__252};
  assign maj__48 = and_60428 ^ a__48 & a__46 ^ and_60345;
  assign temp1__209 = e__49 + S1__52;
  assign ch__52 = e__52 & e__51 ^ ~(e__52 | ~e__50);
  assign value__111 = value__109 + value__110;
  assign s_0__199 = value__69[6:4] ^ value__69[17:15];
  assign s_0__198 = value__69[3:0] ^ value__69[14:11] ^ value__69[31:28];
  assign s_0__197 = value__69[31:21] ^ value__69[10:0] ^ value__69[27:17];
  assign s_0__196 = value__69[20:7] ^ value__69[31:18] ^ value__69[16:3];
  assign s_1__199 = value__108[16:7] ^ value__108[18:9];
  assign s_1__198 = value__108[6:0] ^ value__108[8:2] ^ value__108[31:25];
  assign s_1__197 = value__108[31:30] ^ value__108[1:0] ^ value__108[24:23];
  assign s_1__196 = value__108[29:17] ^ value__108[31:19] ^ value__108[22:10];
  assign temp2__48 = S0__48 + maj__48;
  assign temp1__210 = temp1__209 + ch__52;
  assign temp1__310 = value__111 + 32'h391c_0cb3;
  assign s_0__38 = {s_0__199, s_0__198, s_0__197, s_0__196};
  assign s_1__38 = {s_1__199, s_1__198, s_1__197, s_1__196};
  assign a__49 = temp1__376 + temp2__48;
  assign temp1__212 = temp1__210 + temp1__310;
  assign value__112 = value__66 + s_0__38;
  assign value__113 = value__93 + s_1__38;
  assign e__53 = a__49 + temp1__212;
  assign value__114 = value__112 + value__113;
  assign S0__259 = a__49[1:0] ^ a__49[12:11] ^ a__49[21:20];
  assign S0__258 = a__49[31:21] ^ a__49[10:0] ^ a__49[19:9];
  assign S0__257 = a__49[20:12] ^ a__49[31:23] ^ a__49[8:0];
  assign S0__256 = a__49[11:2] ^ a__49[22:13] ^ a__49[31:22];
  assign and_60498 = a__49 & a__48;
  assign S0__49 = {S0__259, S0__258, S0__257, S0__256};
  assign maj__49 = and_60498 ^ a__49 & a__47 ^ and_60428;
  assign S1__275 = e__53[5:0] ^ e__53[10:5] ^ e__53[24:19];
  assign S1__274 = e__53[31:27] ^ e__53[4:0] ^ e__53[18:14];
  assign S1__273 = e__53[26:13] ^ e__53[31:18] ^ e__53[13:0];
  assign S1__272 = e__53[12:6] ^ e__53[17:11] ^ e__53[31:25];
  assign add_60523 = value__114[31:1] + 31'h276c_5525;
  assign temp2__49 = S0__49 + maj__49;
  assign S1__53 = {S1__275, S1__274, S1__273, S1__272};
  assign ch__53 = e__53 & e__52 ^ ~(e__53 | ~e__51);
  assign temp1__311 = {add_60523, value__114[0]};
  assign a__50 = temp1__373 + temp2__49;
  assign temp1__365 = e__50 + S1__53;
  assign temp1__366 = ch__53 + temp1__311;
  assign temp1__367 = temp1__365 + temp1__366;
  assign S0__263 = a__50[1:0] ^ a__50[12:11] ^ a__50[21:20];
  assign S0__262 = a__50[31:21] ^ a__50[10:0] ^ a__50[19:9];
  assign S0__261 = a__50[20:12] ^ a__50[31:23] ^ a__50[8:0];
  assign S0__260 = a__50[11:2] ^ a__50[22:13] ^ a__50[31:22];
  assign and_60549 = a__50 & a__49;
  assign e__54 = a__50 + temp1__367;
  assign S0__50 = {S0__263, S0__262, S0__261, S0__260};
  assign maj__50 = and_60549 ^ a__50 & a__48 ^ and_60498;
  assign s_0__203 = value__72[6:4] ^ value__72[17:15];
  assign s_0__202 = value__72[3:0] ^ value__72[14:11] ^ value__72[31:28];
  assign s_0__201 = value__72[31:21] ^ value__72[10:0] ^ value__72[27:17];
  assign s_0__200 = value__72[20:7] ^ value__72[31:18] ^ value__72[16:3];
  assign s_1__203 = value__111[16:7] ^ value__111[18:9];
  assign s_1__202 = value__111[6:0] ^ value__111[8:2] ^ value__111[31:25];
  assign s_1__201 = value__111[31:30] ^ value__111[1:0] ^ value__111[24:23];
  assign s_1__200 = value__111[29:17] ^ value__111[31:19] ^ value__111[22:10];
  assign temp2__50 = S0__50 + maj__50;
  assign S1__279 = e__54[5:0] ^ e__54[10:5] ^ e__54[24:19];
  assign S1__278 = e__54[31:27] ^ e__54[4:0] ^ e__54[18:14];
  assign S1__277 = e__54[26:13] ^ e__54[31:18] ^ e__54[13:0];
  assign S1__276 = e__54[12:6] ^ e__54[17:11] ^ e__54[31:25];
  assign s_0__39 = {s_0__203, s_0__202, s_0__201, s_0__200};
  assign s_1__39 = {s_1__203, s_1__202, s_1__201, s_1__200};
  assign a__51 = temp1__370 + temp2__50;
  assign S1__54 = {S1__279, S1__278, S1__277, S1__276};
  assign value__115 = value__69 + s_0__39;
  assign value__116 = value__96 + s_1__39;
  assign temp1__217 = e__51 + S1__54;
  assign ch__54 = e__54 & e__53 ^ ~(e__54 | ~e__52);
  assign value__117 = value__115 + value__116;
  assign S0__267 = a__51[1:0] ^ a__51[12:11] ^ a__51[21:20];
  assign S0__266 = a__51[31:21] ^ a__51[10:0] ^ a__51[19:9];
  assign S0__265 = a__51[20:12] ^ a__51[31:23] ^ a__51[8:0];
  assign S0__264 = a__51[11:2] ^ a__51[22:13] ^ a__51[31:22];
  assign and_60630 = a__51 & a__50;
  assign temp1__218 = temp1__217 + ch__54;
  assign temp1__312 = value__117 + 32'h5b9c_ca4f;
  assign S0__51 = {S0__267, S0__266, S0__265, S0__264};
  assign maj__51 = and_60630 ^ a__51 & a__49 ^ and_60549;
  assign temp1__220 = temp1__218 + temp1__312;
  assign temp2__51 = S0__51 + maj__51;
  assign e__55 = a__51 + temp1__220;
  assign a__52 = temp1__208 + temp2__51;
  assign s_0__207 = value__75[6:4] ^ value__75[17:15];
  assign s_0__206 = value__75[3:0] ^ value__75[14:11] ^ value__75[31:28];
  assign s_0__205 = value__75[31:21] ^ value__75[10:0] ^ value__75[27:17];
  assign s_0__204 = value__75[20:7] ^ value__75[31:18] ^ value__75[16:3];
  assign s_1__207 = value__114[16:7] ^ value__114[18:9];
  assign s_1__206 = value__114[6:0] ^ value__114[8:2] ^ value__114[31:25];
  assign s_1__205 = value__114[31:30] ^ value__114[1:0] ^ value__114[24:23];
  assign s_1__204 = value__114[29:17] ^ value__114[31:19] ^ value__114[22:10];
  assign S1__283 = e__55[5:0] ^ e__55[10:5] ^ e__55[24:19];
  assign S1__282 = e__55[31:27] ^ e__55[4:0] ^ e__55[18:14];
  assign S1__281 = e__55[26:13] ^ e__55[31:18] ^ e__55[13:0];
  assign S1__280 = e__55[12:6] ^ e__55[17:11] ^ e__55[31:25];
  assign s_0__40 = {s_0__207, s_0__206, s_0__205, s_0__204};
  assign s_1__40 = {s_1__207, s_1__206, s_1__205, s_1__204};
  assign S0__271 = a__52[1:0] ^ a__52[12:11] ^ a__52[21:20];
  assign S0__270 = a__52[31:21] ^ a__52[10:0] ^ a__52[19:9];
  assign S0__269 = a__52[20:12] ^ a__52[31:23] ^ a__52[8:0];
  assign S0__268 = a__52[11:2] ^ a__52[22:13] ^ a__52[31:22];
  assign and_60705 = a__52 & a__51;
  assign S1__55 = {S1__283, S1__282, S1__281, S1__280};
  assign value__118 = value__72 + s_0__40;
  assign value__119 = value__99 + s_1__40;
  assign S0__52 = {S0__271, S0__270, S0__269, S0__268};
  assign maj__52 = and_60705 ^ a__52 & a__50 ^ and_60630;
  assign temp1__221 = e__52 + S1__55;
  assign ch__55 = e__55 & e__54 ^ ~(e__55 | ~e__53);
  assign value__120 = value__118 + value__119;
  assign s_0__211 = value__78[6:4] ^ value__78[17:15];
  assign s_0__210 = value__78[3:0] ^ value__78[14:11] ^ value__78[31:28];
  assign s_0__209 = value__78[31:21] ^ value__78[10:0] ^ value__78[27:17];
  assign s_0__208 = value__78[20:7] ^ value__78[31:18] ^ value__78[16:3];
  assign s_1__211 = value__117[16:7] ^ value__117[18:9];
  assign s_1__210 = value__117[6:0] ^ value__117[8:2] ^ value__117[31:25];
  assign s_1__209 = value__117[31:30] ^ value__117[1:0] ^ value__117[24:23];
  assign s_1__208 = value__117[29:17] ^ value__117[31:19] ^ value__117[22:10];
  assign temp2__52 = S0__52 + maj__52;
  assign temp1__222 = temp1__221 + ch__55;
  assign temp1__313 = value__120 + 32'h682e_6ff3;
  assign s_0__41 = {s_0__211, s_0__210, s_0__209, s_0__208};
  assign s_1__41 = {s_1__211, s_1__210, s_1__209, s_1__208};
  assign a__53 = temp1__212 + temp2__52;
  assign temp1__224 = temp1__222 + temp1__313;
  assign value__121 = value__75 + s_0__41;
  assign value__122 = value__102 + s_1__41;
  assign e__56 = a__52 + temp1__224;
  assign value__123 = value__121 + value__122;
  assign S0__275 = a__53[1:0] ^ a__53[12:11] ^ a__53[21:20];
  assign S0__274 = a__53[31:21] ^ a__53[10:0] ^ a__53[19:9];
  assign S0__273 = a__53[20:12] ^ a__53[31:23] ^ a__53[8:0];
  assign S0__272 = a__53[11:2] ^ a__53[22:13] ^ a__53[31:22];
  assign and_60775 = a__53 & a__52;
  assign S0__53 = {S0__275, S0__274, S0__273, S0__272};
  assign maj__53 = and_60775 ^ a__53 & a__51 ^ and_60705;
  assign S1__287 = e__56[5:0] ^ e__56[10:5] ^ e__56[24:19];
  assign S1__286 = e__56[31:27] ^ e__56[4:0] ^ e__56[18:14];
  assign S1__285 = e__56[26:13] ^ e__56[31:18] ^ e__56[13:0];
  assign S1__284 = e__56[12:6] ^ e__56[17:11] ^ e__56[31:25];
  assign add_60800 = value__123[31:1] + 31'h3a47_c177;
  assign temp2__53 = S0__53 + maj__53;
  assign S1__56 = {S1__287, S1__286, S1__285, S1__284};
  assign ch__56 = e__56 & e__55 ^ ~(e__56 | ~e__54);
  assign temp1__314 = {add_60800, value__123[0]};
  assign a__54 = temp1__367 + temp2__53;
  assign temp1__362 = e__53 + S1__56;
  assign temp1__363 = ch__56 + temp1__314;
  assign temp1__364 = temp1__362 + temp1__363;
  assign S0__279 = a__54[1:0] ^ a__54[12:11] ^ a__54[21:20];
  assign S0__278 = a__54[31:21] ^ a__54[10:0] ^ a__54[19:9];
  assign S0__277 = a__54[20:12] ^ a__54[31:23] ^ a__54[8:0];
  assign S0__276 = a__54[11:2] ^ a__54[22:13] ^ a__54[31:22];
  assign and_60826 = a__54 & a__53;
  assign e__57 = a__53 + temp1__364;
  assign S0__54 = {S0__279, S0__278, S0__277, S0__276};
  assign maj__54 = and_60826 ^ a__54 & a__52 ^ and_60775;
  assign s_0__215 = value__81[6:4] ^ value__81[17:15];
  assign s_0__214 = value__81[3:0] ^ value__81[14:11] ^ value__81[31:28];
  assign s_0__213 = value__81[31:21] ^ value__81[10:0] ^ value__81[27:17];
  assign s_0__212 = value__81[20:7] ^ value__81[31:18] ^ value__81[16:3];
  assign s_1__215 = value__120[16:7] ^ value__120[18:9];
  assign s_1__214 = value__120[6:0] ^ value__120[8:2] ^ value__120[31:25];
  assign s_1__213 = value__120[31:30] ^ value__120[1:0] ^ value__120[24:23];
  assign s_1__212 = value__120[29:17] ^ value__120[31:19] ^ value__120[22:10];
  assign temp2__54 = S0__54 + maj__54;
  assign S1__291 = e__57[5:0] ^ e__57[10:5] ^ e__57[24:19];
  assign S1__290 = e__57[31:27] ^ e__57[4:0] ^ e__57[18:14];
  assign S1__289 = e__57[26:13] ^ e__57[31:18] ^ e__57[13:0];
  assign S1__288 = e__57[12:6] ^ e__57[17:11] ^ e__57[31:25];
  assign s_0__42 = {s_0__215, s_0__214, s_0__213, s_0__212};
  assign s_1__42 = {s_1__215, s_1__214, s_1__213, s_1__212};
  assign a__55 = temp1__220 + temp2__54;
  assign S1__57 = {S1__291, S1__290, S1__289, S1__288};
  assign value__124 = value__78 + s_0__42;
  assign value__125 = value__105 + s_1__42;
  assign temp1__229 = e__54 + S1__57;
  assign ch__57 = e__57 & e__56 ^ ~(e__57 | ~e__55);
  assign value__126 = value__124 + value__125;
  assign s_0__219 = value__84[6:4] ^ value__84[17:15];
  assign s_0__218 = value__84[3:0] ^ value__84[14:11] ^ value__84[31:28];
  assign s_0__217 = value__84[31:21] ^ value__84[10:0] ^ value__84[27:17];
  assign s_0__216 = value__84[20:7] ^ value__84[31:18] ^ value__84[16:3];
  assign s_1__219 = value__123[16:7] ^ value__123[18:9];
  assign s_1__218 = value__123[6:0] ^ value__123[8:2] ^ value__123[31:25];
  assign s_1__217 = value__123[31:30] ^ value__123[1:0] ^ value__123[24:23];
  assign s_1__216 = value__123[29:17] ^ value__123[31:19] ^ value__123[22:10];
  assign S0__283 = a__55[1:0] ^ a__55[12:11] ^ a__55[21:20];
  assign S0__282 = a__55[31:21] ^ a__55[10:0] ^ a__55[19:9];
  assign S0__281 = a__55[20:12] ^ a__55[31:23] ^ a__55[8:0];
  assign S0__280 = a__55[11:2] ^ a__55[22:13] ^ a__55[31:22];
  assign and_60936 = a__55 & a__54;
  assign temp1__230 = temp1__229 + ch__57;
  assign temp1__315 = value__126 + 32'h78a5_636f;
  assign s_0__43 = {s_0__219, s_0__218, s_0__217, s_0__216};
  assign s_1__43 = {s_1__219, s_1__218, s_1__217, s_1__216};
  assign S0__55 = {S0__283, S0__282, S0__281, S0__280};
  assign maj__55 = and_60936 ^ a__55 & a__53 ^ and_60826;
  assign temp1__232 = temp1__230 + temp1__315;
  assign value__127 = value__81 + s_0__43;
  assign value__128 = value__108 + s_1__43;
  assign temp2__55 = S0__55 + maj__55;
  assign e__58 = a__54 + temp1__232;
  assign value__129 = value__127 + value__128;
  assign a__56 = temp1__224 + temp2__55;
  assign S1__295 = e__58[5:0] ^ e__58[10:5] ^ e__58[24:19];
  assign S1__294 = e__58[31:27] ^ e__58[4:0] ^ e__58[18:14];
  assign S1__293 = e__58[26:13] ^ e__58[31:18] ^ e__58[13:0];
  assign S1__292 = e__58[12:6] ^ e__58[17:11] ^ e__58[31:25];
  assign add_60984 = value__129[31:2] + 30'h2132_1e05;
  assign S0__287 = a__56[1:0] ^ a__56[12:11] ^ a__56[21:20];
  assign S0__286 = a__56[31:21] ^ a__56[10:0] ^ a__56[19:9];
  assign S0__285 = a__56[20:12] ^ a__56[31:23] ^ a__56[8:0];
  assign S0__284 = a__56[11:2] ^ a__56[22:13] ^ a__56[31:22];
  assign and_61012 = a__56 & a__55;
  assign S1__58 = {S1__295, S1__294, S1__293, S1__292};
  assign ch__58 = e__58 & e__57 ^ ~(e__58 | ~e__56);
  assign temp1__316 = {add_60984, value__129[1:0]};
  assign s_0__223 = value__87[6:4] ^ value__87[17:15];
  assign s_0__222 = value__87[3:0] ^ value__87[14:11] ^ value__87[31:28];
  assign s_0__221 = value__87[31:21] ^ value__87[10:0] ^ value__87[27:17];
  assign s_0__220 = value__87[20:7] ^ value__87[31:18] ^ value__87[16:3];
  assign s_1__223 = value__126[16:7] ^ value__126[18:9];
  assign s_1__222 = value__126[6:0] ^ value__126[8:2] ^ value__126[31:25];
  assign s_1__221 = value__126[31:30] ^ value__126[1:0] ^ value__126[24:23];
  assign s_1__220 = value__126[29:17] ^ value__126[31:19] ^ value__126[22:10];
  assign S0__56 = {S0__287, S0__286, S0__285, S0__284};
  assign maj__56 = and_61012 ^ a__56 & a__54 ^ and_60936;
  assign temp1__359 = e__55 + S1__58;
  assign temp1__360 = ch__58 + temp1__316;
  assign s_0__44 = {s_0__223, s_0__222, s_0__221, s_0__220};
  assign s_1__44 = {s_1__223, s_1__222, s_1__221, s_1__220};
  assign temp2__56 = S0__56 + maj__56;
  assign temp1__361 = temp1__359 + temp1__360;
  assign value__130 = value__84 + s_0__44;
  assign value__131 = value__111 + s_1__44;
  assign a__57 = temp1__364 + temp2__56;
  assign e__59 = a__55 + temp1__361;
  assign value__132 = value__130 + value__131;
  assign S0__291 = a__57[1:0] ^ a__57[12:11] ^ a__57[21:20];
  assign S0__290 = a__57[31:21] ^ a__57[10:0] ^ a__57[19:9];
  assign S0__289 = a__57[20:12] ^ a__57[31:23] ^ a__57[8:0];
  assign S0__288 = a__57[11:2] ^ a__57[22:13] ^ a__57[31:22];
  assign and_61069 = a__57 & a__56;
  assign S1__299 = e__59[5:0] ^ e__59[10:5] ^ e__59[24:19];
  assign S1__298 = e__59[31:27] ^ e__59[4:0] ^ e__59[18:14];
  assign S1__297 = e__59[26:13] ^ e__59[31:18] ^ e__59[13:0];
  assign S1__296 = e__59[12:6] ^ e__59[17:11] ^ e__59[31:25];
  assign add_61077 = value__132[31:3] + 29'h1198_e041;
  assign S0__57 = {S0__291, S0__290, S0__289, S0__288};
  assign maj__57 = and_61069 ^ a__57 & a__55 ^ and_61012;
  assign S1__59 = {S1__299, S1__298, S1__297, S1__296};
  assign ch__59 = e__59 & e__58 ^ ~(e__59 | ~e__57);
  assign temp1__317 = {add_61077, value__132[2:0]};
  assign s_0__227 = value__90[6:4] ^ value__90[17:15];
  assign s_0__226 = value__90[3:0] ^ value__90[14:11] ^ value__90[31:28];
  assign s_0__225 = value__90[31:21] ^ value__90[10:0] ^ value__90[27:17];
  assign s_0__224 = value__90[20:7] ^ value__90[31:18] ^ value__90[16:3];
  assign s_1__227 = value__129[16:7] ^ value__129[18:9];
  assign s_1__226 = value__129[6:0] ^ value__129[8:2] ^ value__129[31:25];
  assign s_1__225 = value__129[31:30] ^ value__129[1:0] ^ value__129[24:23];
  assign s_1__224 = value__129[29:17] ^ value__129[31:19] ^ value__129[22:10];
  assign temp2__57 = S0__57 + maj__57;
  assign temp1__356 = e__56 + S1__59;
  assign temp1__357 = ch__59 + temp1__317;
  assign s_0__45 = {s_0__227, s_0__226, s_0__225, s_0__224};
  assign s_1__45 = {s_1__227, s_1__226, s_1__225, s_1__224};
  assign a__58 = temp1__232 + temp2__57;
  assign temp1__358 = temp1__356 + temp1__357;
  assign value__133 = value__87 + s_0__45;
  assign value__134 = value__114 + s_1__45;
  assign e__60 = a__56 + temp1__358;
  assign value__135 = value__133 + value__134;
  assign S0__295 = a__58[1:0] ^ a__58[12:11] ^ a__58[21:20];
  assign S0__294 = a__58[31:21] ^ a__58[10:0] ^ a__58[19:9];
  assign S0__293 = a__58[20:12] ^ a__58[31:23] ^ a__58[8:0];
  assign S0__292 = a__58[11:2] ^ a__58[22:13] ^ a__58[31:22];
  assign and_61140 = a__58 & a__57;
  assign S0__58 = {S0__295, S0__294, S0__293, S0__292};
  assign maj__58 = and_61140 ^ a__58 & a__56 ^ and_61069;
  assign S1__303 = e__60[5:0] ^ e__60[10:5] ^ e__60[24:19];
  assign S1__302 = e__60[31:27] ^ e__60[4:0] ^ e__60[18:14];
  assign S1__301 = e__60[26:13] ^ e__60[31:18] ^ e__60[13:0];
  assign S1__300 = e__60[12:6] ^ e__60[17:11] ^ e__60[31:25];
  assign add_61165 = value__135[31:1] + 31'h485f_7ffd;
  assign temp2__58 = S0__58 + maj__58;
  assign S1__60 = {S1__303, S1__302, S1__301, S1__300};
  assign ch__60 = e__60 & e__59 ^ ~(e__60 | ~e__58);
  assign temp1__318 = {add_61165, value__135[0]};
  assign a__59 = temp1__361 + temp2__58;
  assign temp1__353 = e__57 + S1__60;
  assign temp1__354 = ch__60 + temp1__318;
  assign temp1__355 = temp1__353 + temp1__354;
  assign S0__299 = a__59[1:0] ^ a__59[12:11] ^ a__59[21:20];
  assign S0__298 = a__59[31:21] ^ a__59[10:0] ^ a__59[19:9];
  assign S0__297 = a__59[20:12] ^ a__59[31:23] ^ a__59[8:0];
  assign S0__296 = a__59[11:2] ^ a__59[22:13] ^ a__59[31:22];
  assign and_61191 = a__59 & a__58;
  assign e__61 = a__57 + temp1__355;
  assign S0__59 = {S0__299, S0__298, S0__297, S0__296};
  assign maj__59 = and_61191 ^ a__59 & a__57 ^ and_61140;
  assign s_0__231 = value__93[6:4] ^ value__93[17:15];
  assign s_0__230 = value__93[3:0] ^ value__93[14:11] ^ value__93[31:28];
  assign s_0__229 = value__93[31:21] ^ value__93[10:0] ^ value__93[27:17];
  assign s_0__228 = value__93[20:7] ^ value__93[31:18] ^ value__93[16:3];
  assign s_1__231 = value__132[16:7] ^ value__132[18:9];
  assign s_1__230 = value__132[6:0] ^ value__132[8:2] ^ value__132[31:25];
  assign s_1__229 = value__132[31:30] ^ value__132[1:0] ^ value__132[24:23];
  assign s_1__228 = value__132[29:17] ^ value__132[31:19] ^ value__132[22:10];
  assign temp2__59 = S0__59 + maj__59;
  assign S1__307 = e__61[5:0] ^ e__61[10:5] ^ e__61[24:19];
  assign S1__306 = e__61[31:27] ^ e__61[4:0] ^ e__61[18:14];
  assign S1__305 = e__61[26:13] ^ e__61[31:18] ^ e__61[13:0];
  assign S1__304 = e__61[12:6] ^ e__61[17:11] ^ e__61[31:25];
  assign s_0__46 = {s_0__231, s_0__230, s_0__229, s_0__228};
  assign s_1__46 = {s_1__231, s_1__230, s_1__229, s_1__228};
  assign a__60 = temp1__358 + temp2__59;
  assign S1__61 = {S1__307, S1__306, S1__305, S1__304};
  assign value__136 = value__90 + s_0__46;
  assign value__137 = value__117 + s_1__46;
  assign temp1__245 = e__58 + S1__61;
  assign ch__61 = e__61 & e__60 ^ ~(e__61 | ~e__59);
  assign value__138 = value__136 + value__137;
  assign S0__303 = a__60[1:0] ^ a__60[12:11] ^ a__60[21:20];
  assign S0__302 = a__60[31:21] ^ a__60[10:0] ^ a__60[19:9];
  assign S0__301 = a__60[20:12] ^ a__60[31:23] ^ a__60[8:0];
  assign S0__300 = a__60[11:2] ^ a__60[22:13] ^ a__60[31:22];
  assign and_61272 = a__60 & a__59;
  assign temp1__246 = temp1__245 + ch__61;
  assign temp1__319 = value__138 + 32'ha450_6ceb;
  assign S0__60 = {S0__303, S0__302, S0__301, S0__300};
  assign maj__60 = and_61272 ^ a__60 & a__58 ^ and_61191;
  assign temp1__248 = temp1__246 + temp1__319;
  assign temp2__60 = S0__60 + maj__60;
  assign e__62 = a__58 + temp1__248;
  assign a__61 = temp1__355 + temp2__60;
  assign S1__311 = e__62[5:0] ^ e__62[10:5] ^ e__62[24:19];
  assign S1__310 = e__62[31:27] ^ e__62[4:0] ^ e__62[18:14];
  assign S1__309 = e__62[26:13] ^ e__62[31:18] ^ e__62[13:0];
  assign S1__308 = e__62[12:6] ^ e__62[17:11] ^ e__62[31:25];
  assign s_0__235 = value__96[6:4] ^ value__96[17:15];
  assign s_0__234 = value__96[3:0] ^ value__96[14:11] ^ value__96[31:28];
  assign s_0__233 = value__96[31:21] ^ value__96[10:0] ^ value__96[27:17];
  assign s_0__232 = value__96[20:7] ^ value__96[31:18] ^ value__96[16:3];
  assign s_1__235 = value__135[16:7] ^ value__135[18:9];
  assign s_1__234 = value__135[6:0] ^ value__135[8:2] ^ value__135[31:25];
  assign s_1__233 = value__135[31:30] ^ value__135[1:0] ^ value__135[24:23];
  assign s_1__232 = value__135[29:17] ^ value__135[31:19] ^ value__135[22:10];
  assign S0__307 = a__61[1:0] ^ a__61[12:11] ^ a__61[21:20];
  assign S0__306 = a__61[31:21] ^ a__61[10:0] ^ a__61[19:9];
  assign S0__305 = a__61[20:12] ^ a__61[31:23] ^ a__61[8:0];
  assign S0__304 = a__61[11:2] ^ a__61[22:13] ^ a__61[31:22];
  assign and_61346 = a__61 & a__60;
  assign S1__62 = {S1__311, S1__310, S1__309, S1__308};
  assign ch__62 = e__62 & e__61 ^ ~(e__62 | ~e__60);
  assign s_0__47 = {s_0__235, s_0__234, s_0__233, s_0__232};
  assign s_1__47 = {s_1__235, s_1__234, s_1__233, s_1__232};
  assign S0__61 = {S0__307, S0__306, S0__305, S0__304};
  assign maj__61 = and_61346 ^ a__61 & a__59 ^ and_61272;
  assign temp1__346 = e__59 + S1__62;
  assign temp1__347 = ch__62 + value__93;
  assign temp1__348 = s_0__47 + value__120;
  assign temp1__349 = s_1__47 + 32'hbef9_a3f7;
  assign temp2__61 = S0__61 + maj__61;
  assign temp1__350 = temp1__346 + temp1__347;
  assign temp1__351 = temp1__348 + temp1__349;
  assign a__62 = temp1__248 + temp2__61;
  assign temp1__352 = temp1__350 + temp1__351;
  assign e__63 = a__59 + temp1__352;
  assign s_1__236 = value__138[29:17] ^ value__138[31:19] ^ value__138[22:10];
  assign S0__311 = a__62[1:0] ^ a__62[12:11] ^ a__62[21:20];
  assign S0__310 = a__62[31:21] ^ a__62[10:0] ^ a__62[19:9];
  assign S0__309 = a__62[20:12] ^ a__62[31:23] ^ a__62[8:0];
  assign S0__308 = a__62[11:2] ^ a__62[22:13] ^ a__62[31:22];
  assign and_61393 = a__62 & a__61;
  assign s_1__239 = value__138[16:7] ^ value__138[18:9];
  assign s_1__238 = value__138[6:0] ^ value__138[8:2] ^ value__138[31:25];
  assign s_1__237 = value__138[31:30] ^ value__138[1:0] ^ value__138[24:23];
  assign S0__62 = {S0__311, S0__310, S0__309, S0__308};
  assign maj__62 = and_61393 ^ a__62 & a__60 ^ and_61346;
  assign S1__315 = e__63[5:0] ^ e__63[10:5] ^ e__63[24:19];
  assign S1__314 = e__63[31:27] ^ e__63[4:0] ^ e__63[18:14];
  assign S1__313 = e__63[26:13] ^ e__63[31:18] ^ e__63[13:0];
  assign S1__312 = e__63[12:6] ^ e__63[17:11] ^ e__63[31:25];
  assign s_0__239 = value__99[6:4] ^ value__99[17:15];
  assign s_0__238 = value__99[3:0] ^ value__99[14:11] ^ value__99[31:28];
  assign s_0__237 = value__99[31:21] ^ value__99[10:0] ^ value__99[27:17];
  assign s_0__236 = value__99[20:7] ^ value__99[31:18] ^ value__99[16:3];
  assign temp2__62 = S0__62 + maj__62;
  assign S1__63 = {S1__315, S1__314, S1__313, S1__312};
  assign ch__63 = e__63 & e__62 ^ ~(e__63 | ~e__61);
  assign s_0__240 = {s_0__239, s_0__238, s_0__237, s_0__236};
  assign add_61441 = {s_1__239, s_1__238, s_1__237, s_1__236[12:1]} + 31'h6338_bc79;
  assign a__63 = temp1__352 + temp2__62;
  assign temp1__339 = e__60 + S1__63;
  assign temp1__340 = ch__63 + value__96;
  assign temp1__341 = s_0__240 + value__123;
  assign temp1__342 = {add_61441, s_1__236[0]};
  assign temp1__343 = temp1__339 + temp1__340;
  assign temp1__344 = temp1__341 + temp1__342;
  assign S0__315 = a__63[1:0] ^ a__63[12:11] ^ a__63[21:20];
  assign S0__314 = a__63[31:21] ^ a__63[10:0] ^ a__63[19:9];
  assign S0__313 = a__63[20:12] ^ a__63[31:23] ^ a__63[8:0];
  assign S0__312 = a__63[11:2] ^ a__63[22:13] ^ a__63[31:22];
  assign temp1__345 = temp1__343 + temp1__344;
  assign S0__63 = {S0__315, S0__314, S0__313, S0__312};
  assign maj__63 = a__63 & a__62 ^ a__63 & a__61 ^ and_61393;
  assign b__68 = 32'h6a09_e667;
  assign add_61478 = temp1__345 + S0__63;
  assign add_61479 = maj__63 + b__68;
  assign c__66 = 32'hbb67_ae85;
  assign add_61481 = a__62[31:1] + 31'h1e37_79b9;
  assign add_61483 = a__61[31:1] + 31'h52a7_fa9d;
  assign e__64 = a__60 + temp1__345;
  assign f__66 = 32'h510e_527f;
  assign add_61487 = e__63[31:2] + 30'h26c1_5a23;
  assign h__1 = 32'h1f83_d9ab;
  assign h7 = 32'h5be0_cd19;
  assign add_61491 = add_61478 + add_61479;
  assign add_61492 = a__63 + c__66;
  assign add_61495 = e__64 + f__66;
  assign add_61497 = e__62 + h__1;
  assign add_61498 = e__61 + h7;
  assign out = {add_61491, add_61492, {add_61481, a__62[0]}, {add_61483, a__61[0]}, add_61495, {add_61487, e__63[1:0]}, add_61497, add_61498};
endmodule
