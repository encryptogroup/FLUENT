module __f32add__main(
  input wire [31:0] x,
  input wire [31:0] y,
  output wire [31:0] out
);
  wire [22:0] x_fraction__1;
  wire [7:0] x_bexp__1;
  wire [22:0] y_fraction__3;
  wire [7:0] y_bexp__1;
  wire [5:0] add_1786;
  wire ugt_1788;
  wire [5:0] add_1792;
  wire [27:0] wide_x;
  wire [7:0] greater_exp_bexp;
  wire [27:0] wide_y;
  wire [27:0] wide_x__1;
  wire [7:0] sub_1802;
  wire [27:0] wide_y__1;
  wire [7:0] sub_1804;
  wire [27:0] dropped_x;
  wire [27:0] dropped_y;
  wire [7:0] shift_x;
  wire sticky_x;
  wire [7:0] shift_y;
  wire sticky_y;
  wire y_sign__1;
  wire x_sign__1;
  wire [27:0] shifted_x;
  wire [27:0] shifted_y;
  wire greater_exp_sign;
  wire [27:0] addend_x;
  wire [27:0] addend_y;
  wire [27:0] addend_x__1;
  wire [27:0] addend_y__1;
  wire [28:0] fraction;
  wire [27:0] abs_fraction;
  wire [27:0] reverse_1839;
  wire [28:0] one_hot_1840;
  wire [4:0] encode_1841;
  wire carry_bit;
  wire cancel;
  wire and_1850;
  wire and_1851;
  wire and_1852;
  wire [27:0] leading_zeroes;
  wire [26:0] carry_fraction;
  wire [27:0] add_1865;
  wire [3:0] concat_1866;
  wire [26:0] carry_fraction__1;
  wire [26:0] cancel_fraction;
  wire [26:0] shifted_fraction;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [24:0] add_1882;
  wire do_round_up;
  wire [27:0] rounded_fraction;
  wire rounding_carry;
  wire [8:0] add_1893;
  wire [9:0] add_1898;
  wire [9:0] wide_exponent;
  wire [9:0] wide_exponent__1;
  wire [7:0] max_exp__3;
  wire [7:0] max_exp__4;
  wire [7:0] max_exp__1;
  wire [7:0] max_exp__2;
  wire [8:0] wide_exponent__2;
  wire ne_1918;
  wire ne_1920;
  wire eq_1921;
  wire eq_1922;
  wire eq_1923;
  wire eq_1924;
  wire has_pos_inf;
  wire has_neg_inf;
  wire fraction_is_zero;
  wire [2:0] add_1949;
  wire and_1951;
  wire and_1952;
  wire nor_1958;
  wire [27:0] shrl_1959;
  wire is_result_nan;
  wire is_operand_inf;
  wire result_sign;
  wire [22:0] result_fraction;
  wire result_sign__1;
  wire [7:0] max_exp__5;
  wire [22:0] result_fraction__3;
  wire [22:0] fraction_high_bit;
  wire result_sign__3;
  wire [7:0] result_exponent__2;
  wire [22:0] result_fraction__4;
  assign x_fraction__1 = x[22:0];
  assign x_bexp__1 = x[30:23];
  assign y_fraction__3 = y[22:0];
  assign y_bexp__1 = y[30:23];
  assign add_1786 = x_bexp__1[7:2] + 6'h07;
  assign ugt_1788 = x_bexp__1 > y_bexp__1;
  assign add_1792 = y_bexp__1[7:2] + 6'h07;
  assign wide_x = {{2'h0, x_fraction__1} | 25'h080_0000, 3'h0};
  assign greater_exp_bexp = ugt_1788 ? x_bexp__1 : y_bexp__1;
  assign wide_y = {{2'h0, y_fraction__3} | 25'h080_0000, 3'h0};
  assign wide_x__1 = wide_x & {28{x_bexp__1 != 8'h00}};
  assign sub_1802 = {add_1786, x_bexp__1[1:0]} - greater_exp_bexp;
  assign wide_y__1 = wide_y & {28{y_bexp__1 != 8'h00}};
  assign sub_1804 = {add_1792, y_bexp__1[1:0]} - greater_exp_bexp;
  assign dropped_x = sub_1802 >= 8'h1c ? 28'h000_0000 : wide_x__1 << sub_1802;
  assign dropped_y = sub_1804 >= 8'h1c ? 28'h000_0000 : wide_y__1 << sub_1804;
  assign shift_x = greater_exp_bexp - x_bexp__1;
  assign sticky_x = dropped_x[27:3] != 25'h000_0000;
  assign shift_y = greater_exp_bexp - y_bexp__1;
  assign sticky_y = dropped_y[27:3] != 25'h000_0000;
  assign y_sign__1 = y[31:31];
  assign x_sign__1 = x[31:31];
  assign shifted_x = shift_x >= 8'h1c ? 28'h000_0000 : wide_x__1 >> shift_x;
  assign shifted_y = shift_y >= 8'h1c ? 28'h000_0000 : wide_y__1 >> shift_y;
  assign greater_exp_sign = ugt_1788 ? x_sign__1 : y_sign__1;
  assign addend_x = shifted_x | {27'h000_0000, sticky_x};
  assign addend_y = shifted_y | {27'h000_0000, sticky_y};
  assign addend_x__1 = x_sign__1 ^ greater_exp_sign ? -addend_x : addend_x;
  assign addend_y__1 = y_sign__1 ^ greater_exp_sign ? -addend_y : addend_y;
  assign fraction = {{1{addend_x__1[27]}}, addend_x__1} + {{1{addend_y__1[27]}}, addend_y__1};
  assign abs_fraction = fraction[28] ? -fraction[27:0] : fraction[27:0];
  assign reverse_1839 = {abs_fraction[0], abs_fraction[1], abs_fraction[2], abs_fraction[3], abs_fraction[4], abs_fraction[5], abs_fraction[6], abs_fraction[7], abs_fraction[8], abs_fraction[9], abs_fraction[10], abs_fraction[11], abs_fraction[12], abs_fraction[13], abs_fraction[14], abs_fraction[15], abs_fraction[16], abs_fraction[17], abs_fraction[18], abs_fraction[19], abs_fraction[20], abs_fraction[21], abs_fraction[22], abs_fraction[23], abs_fraction[24], abs_fraction[25], abs_fraction[26], abs_fraction[27]};
  assign one_hot_1840 = {reverse_1839[27:0] == 28'h000_0000, reverse_1839[27] && reverse_1839[26:0] == 27'h000_0000, reverse_1839[26] && reverse_1839[25:0] == 26'h000_0000, reverse_1839[25] && reverse_1839[24:0] == 25'h000_0000, reverse_1839[24] && reverse_1839[23:0] == 24'h00_0000, reverse_1839[23] && reverse_1839[22:0] == 23'h00_0000, reverse_1839[22] && reverse_1839[21:0] == 22'h00_0000, reverse_1839[21] && reverse_1839[20:0] == 21'h00_0000, reverse_1839[20] && reverse_1839[19:0] == 20'h0_0000, reverse_1839[19] && reverse_1839[18:0] == 19'h0_0000, reverse_1839[18] && reverse_1839[17:0] == 18'h0_0000, reverse_1839[17] && reverse_1839[16:0] == 17'h0_0000, reverse_1839[16] && reverse_1839[15:0] == 16'h0000, reverse_1839[15] && reverse_1839[14:0] == 15'h0000, reverse_1839[14] && reverse_1839[13:0] == 14'h0000, reverse_1839[13] && reverse_1839[12:0] == 13'h0000, reverse_1839[12] && reverse_1839[11:0] == 12'h000, reverse_1839[11] && reverse_1839[10:0] == 11'h000, reverse_1839[10] && reverse_1839[9:0] == 10'h000, reverse_1839[9] && reverse_1839[8:0] == 9'h000, reverse_1839[8] && reverse_1839[7:0] == 8'h00, reverse_1839[7] && reverse_1839[6:0] == 7'h00, reverse_1839[6] && reverse_1839[5:0] == 6'h00, reverse_1839[5] && reverse_1839[4:0] == 5'h00, reverse_1839[4] && reverse_1839[3:0] == 4'h0, reverse_1839[3] && reverse_1839[2:0] == 3'h0, reverse_1839[2] && reverse_1839[1:0] == 2'h0, reverse_1839[1] && !reverse_1839[0], reverse_1839[0]};
  assign encode_1841 = {one_hot_1840[16] | one_hot_1840[17] | one_hot_1840[18] | one_hot_1840[19] | one_hot_1840[20] | one_hot_1840[21] | one_hot_1840[22] | one_hot_1840[23] | one_hot_1840[24] | one_hot_1840[25] | one_hot_1840[26] | one_hot_1840[27] | one_hot_1840[28], one_hot_1840[8] | one_hot_1840[9] | one_hot_1840[10] | one_hot_1840[11] | one_hot_1840[12] | one_hot_1840[13] | one_hot_1840[14] | one_hot_1840[15] | one_hot_1840[24] | one_hot_1840[25] | one_hot_1840[26] | one_hot_1840[27] | one_hot_1840[28], one_hot_1840[4] | one_hot_1840[5] | one_hot_1840[6] | one_hot_1840[7] | one_hot_1840[12] | one_hot_1840[13] | one_hot_1840[14] | one_hot_1840[15] | one_hot_1840[20] | one_hot_1840[21] | one_hot_1840[22] | one_hot_1840[23] | one_hot_1840[28], one_hot_1840[2] | one_hot_1840[3] | one_hot_1840[6] | one_hot_1840[7] | one_hot_1840[10] | one_hot_1840[11] | one_hot_1840[14] | one_hot_1840[15] | one_hot_1840[18] | one_hot_1840[19] | one_hot_1840[22] | one_hot_1840[23] | one_hot_1840[26] | one_hot_1840[27], one_hot_1840[1] | one_hot_1840[3] | one_hot_1840[5] | one_hot_1840[7] | one_hot_1840[9] | one_hot_1840[11] | one_hot_1840[13] | one_hot_1840[15] | one_hot_1840[17] | one_hot_1840[19] | one_hot_1840[21] | one_hot_1840[23] | one_hot_1840[25] | one_hot_1840[27]};
  assign carry_bit = abs_fraction[27];
  assign cancel = encode_1841[1] | encode_1841[2] | encode_1841[3] | encode_1841[4];
  assign and_1850 = ~carry_bit & ~cancel;
  assign and_1851 = ~carry_bit & cancel;
  assign and_1852 = carry_bit & ~cancel;
  assign leading_zeroes = {23'h00_0000, encode_1841};
  assign carry_fraction = abs_fraction[27:1];
  assign add_1865 = leading_zeroes + 28'hfff_ffff;
  assign concat_1866 = {~and_1850 & ~and_1851 & ~and_1852, and_1850, and_1851, and_1852};
  assign carry_fraction__1 = carry_fraction | {26'h000_0000, abs_fraction[0]};
  assign cancel_fraction = add_1865 >= 28'h000_001b ? 27'h000_0000 : abs_fraction[26:0] << add_1865;
  assign shifted_fraction = carry_fraction__1 & {27{concat_1866[0]}} | cancel_fraction & {27{concat_1866[1]}} | abs_fraction[26:0] & {27{concat_1866[2]}} | 27'h000_029a & {27{concat_1866[3]}};
  assign normal_chunk = shifted_fraction[2:0];
  assign half_way_chunk = shifted_fraction[3:2];
  assign add_1882 = {1'h0, shifted_fraction[26:3]} + 25'h000_0001;
  assign do_round_up = normal_chunk > 3'h4 | half_way_chunk == 2'h3;
  assign rounded_fraction = do_round_up ? {add_1882, normal_chunk} : {1'h0, shifted_fraction};
  assign rounding_carry = rounded_fraction[27];
  assign add_1893 = {1'h0, greater_exp_bexp} + {8'h00, rounding_carry};
  assign add_1898 = {1'h0, add_1893} + 10'h001;
  assign wide_exponent = add_1898 - {5'h00, encode_1841};
  assign wide_exponent__1 = wide_exponent & {10{fraction != 29'h0000_0000}};
  assign max_exp__3 = 8'hff;
  assign max_exp__4 = 8'hff;
  assign max_exp__1 = 8'hff;
  assign max_exp__2 = 8'hff;
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign ne_1918 = x_fraction__1 != 23'h00_0000;
  assign ne_1920 = y_fraction__3 != 23'h00_0000;
  assign eq_1921 = x_bexp__1 == max_exp__1;
  assign eq_1922 = x_fraction__1 == 23'h00_0000;
  assign eq_1923 = y_bexp__1 == max_exp__2;
  assign eq_1924 = y_fraction__3 == 23'h00_0000;
  assign has_pos_inf = ~(x_bexp__1 != max_exp__3 | ne_1918 | x_sign__1) | ~(y_bexp__1 != max_exp__4 | ne_1920 | y_sign__1);
  assign has_neg_inf = eq_1921 & eq_1922 & x_sign__1 | eq_1923 & eq_1924 & y_sign__1;
  assign fraction_is_zero = fraction == 29'h0000_0000;
  assign add_1949 = {2'h0, rounding_carry} + 3'h3;
  assign and_1951 = eq_1921 & eq_1922;
  assign and_1952 = eq_1923 & eq_1924;
  assign nor_1958 = ~(wide_exponent__2[8] | wide_exponent__2[0] & wide_exponent__2[1] & wide_exponent__2[2] & wide_exponent__2[3] & wide_exponent__2[4] & wide_exponent__2[5] & wide_exponent__2[6] & wide_exponent__2[7]);
  assign shrl_1959 = rounded_fraction >> add_1949;
  assign is_result_nan = eq_1921 & ne_1918 | eq_1923 & ne_1920 | has_pos_inf & has_neg_inf;
  assign is_operand_inf = and_1951 | and_1952;
  assign result_sign = ~(~fraction[28] | greater_exp_sign) | ~(fraction[28] | fraction_is_zero | ~greater_exp_sign);
  assign result_fraction = shrl_1959[22:0];
  assign result_sign__1 = is_operand_inf ? ~has_pos_inf : result_sign;
  assign max_exp__5 = 8'hff;
  assign result_fraction__3 = result_fraction & {23{~(~(wide_exponent__2[1] | wide_exponent__2[2] | wide_exponent__2[3] | wide_exponent__2[4] | wide_exponent__2[5] | wide_exponent__2[6] | wide_exponent__2[7] | wide_exponent__2[8] | wide_exponent__2[0]))}} & {23{nor_1958}} & {23{~(and_1951 | and_1952)}};
  assign fraction_high_bit = 23'h40_0000;
  assign result_sign__3 = ~is_result_nan & result_sign__1;
  assign result_exponent__2 = is_result_nan | is_operand_inf | ~nor_1958 ? max_exp__5 : wide_exponent__2[7:0];
  assign result_fraction__4 = is_result_nan ? fraction_high_bit : result_fraction__3;
  assign out = {result_sign__3, result_exponent__2, result_fraction__4};
endmodule
